  X � 
   % 0� 
   % 0 LIB  >A�7KƧ�9D�/��ZT � 
   % 0� 
   % 0 $$$CONTEXT_INFO$$$ 
  res_poly$4          +  ,PCELL=res_poly +  ,P(w)=##0.35  +  ,,P(type)='sky130_fd_pr__res_high_po_0p35' +  ,P(res_value)=##784.99925 +  ,P(len)=##0.25  +  ,P(gr)=false  +  ,P(area)=##0.0875 +   ,LIB=skywater130    
  res_poly$3          +  ,PCELL=res_poly +  ,P(w)=##0.35  +  ,,P(type)='sky130_fd_pr__res_high_po_0p35' +  ,P(res_value)=##1569.9985 +  ,P(len)=##0.5 +  ,P(gr)=false  +  ,P(area)=##0.175  +   ,LIB=skywater130    
  
pfet$6          +  ,PCELL=pfet +  ,P(w)=##40  +  &,P(type)='sky130_fd_pr__pfet_01v8'  +  ,P(sd_con_col)=#l3  +  ,P(perim)=##88  + 
 ,P(patt)='' + 	 ,P(nf)=#l1  +  ,P(l)=##4 +  ,P(interdig)=true +  ,P(inter_sd_l)=##0.5  +  ,P(grw)=##0.17  +  ,P(gate_con_pos)='top'  +  ,P(con_bet_fin)=true  +  ,P(bulk)='bulk tie' +  ,P(area)=##160  +   ,LIB=skywater130    
  nfet$10           +  ,PCELL=nfet +  ,P(w)=##30  +  &,P(type)='sky130_fd_pr__nfet_01v8'  +  ,P(sd_con_col)=##2  +  ,P(perim)=##64  + 
 ,P(patt)='' + 	 ,P(nf)=#l1  +  ,P(l)=##2 +  ,P(interdig)=true +  ,P(inter_sd_l)=##0.5  +  ,P(grw)=##0.3 +  ,P(gate_con_pos)='top'  +  ,P(con_bet_fin)=true  +  ,P(bulk)='None' +  ,P(area)=##60 +   ,LIB=skywater130    
  nfet          +  ,PCELL=nfet +  ,P(w)=##1 +  &,P(type)='sky130_fd_pr__nfet_01v8'  +  ,P(sd_con_col)=##1  +  ,P(perim)=##2.4 + 
 ,P(patt)='' + 	 ,P(nf)=#l1  +  ,P(l)=##0.2 +  ,P(interdig)=true +  ,P(inter_sd_l)=##0.5  +  ,P(grw)=##0.3 +  ,P(gate_con_pos)='top'  +  ,P(con_bet_fin)=true  +  ,P(bulk)='bulk tie' +  ,P(area)=##0.2  +   ,LIB=skywater130      � 
   % 0� 
   % 0 res_poly$4    B   ,���Q������Q  �   �  �   �������Q���      D   ,����   �����  �   }  �   }   �����   �      D   ,�������1�������i   }���i   }���1�������1      _   ,������������  	L    	L  ������������      C   ,���Q   }���Q  �   �  �   �   }���Q   }      C   ,���Q������Q����   �����   �������Q���      ^   ,������������  	[    	[  ������������      C  , ,����   �����  �   U  �   U   �����   �      C  , ,����  D����  �   U  �   U  D����  D      C  , ,����  �����  V   U  V   U  �����  �      C  , ,����  ����  �   U  �   U  ����        C  , ,����  |����  &   U  &   U  |����  |      C  , ,����  �����  �   U  �   U  �����  �      C  , ,�������w�������!   U���!   U���w�������w      C  , ,����������������   U����   U������������      C  , ,�������G��������   U����   U���G�������G      C  , ,���������������Y   U���Y   U������������      C  , ,���������������   U����   U����������      C  , ,��������������)   U���)   U����������      B  , ,����   �����  �   _  �   _   �����   �      B  , ,�������c�������3   _���3   _���c�������c      B   ,���Q���G���Q   �   �   �   ����G���Q���G      V   ,�������K����  	�  {  	�  {���K�������K     � 
   % 0� 
   % 0 res_poly$3    B   ,���Q�������Q  	j   �  	j   ��������Q����      D   ,����  ����  	L   }  	L   }  ����        D   ,����������������   }����   }������������      _   ,�������7����  	�    	�  ���7�������7      C   ,���Q   ����Q  	j   �  	j   �   ����Q   �      C   ,���Q�������Q���   ����   ��������Q����      ^   ,�������(����  	�    	�  ���(�������(      C  , ,����  Y����     U     U  Y����  Y      C  , ,����  �����  k   U  k   U  �����  �      C  , ,����  )����  �   U  �   U  )����  )      C  , ,����  �����  ;   U  ;   U  �����  �      C  , ,����  �����  �   U  �   U  �����  �      C  , ,����  a����  	   U  	   U  a����  a      C  , ,����������������   U����   U������������      C  , ,�������b�������   U���   U���b�������b      C  , ,���������������t   U���t   U������������      C  , ,�������2��������   U����   U���2�������2      C  , ,���������������D   U���D   U������������      C  , ,���������������   U����   U����������      B  , ,����  J����  	   _  	   _  J����  J      B  , ,����������������   _����   _������������      B   ,���Q�������Q  6   �  6   ��������Q����      V   ,������������  
2  {  
2  {������������     � 
   % 0� 
   % 0 sky130_fd_sc_hd__buf_16     B  l  �   i  �  
7  !  
7  !    /    /  
7  �  
7  �    �    �  
7  i  
7  i    w    w  
7    
7            
7  �  
7  �    	�    	�  
7  
U  
7  
U   i  	�   i  	�    �    �   i     i             i  w   i  w    i    i   i  �   i  �    �    �   i  /   i  /    !    !   i  �   i      B    c   i  c  
7  �  
7  �          
7  �  
7  �    �    �  
7  A  
7  A    O    O  
7  �  
7  �    �    �  
7  �  
7  �    �    �  
7  -  
7  -    ;    ;  
7  �  
7  �    �    �  
7  u  
7  u    �    �  
7    
7      '    '  
7  �  
7  �    �    �  
7  a  
7  a    o    o  
7    
7            
7  �  
7  �     �     �  
7  !M  
7  !M    "[    "[  
7  "�  
7  "�    #�    #�  
7  $�  
7  $�    $�    $�    $�    $�   i  #�   i  #�    "�    "�   i  "[   i  "[    !M    !M   i   �   i   �    �    �   i     i             i  o   i  o    a    a   i  �   i  �    �    �   i  '   i  '           i  �   i  �    u    u   i  �   i  �    �    �   i  ;   i  ;    -    -   i  �   i  �    �    �   i  �   i  �    �    �   i  O   i  O    A    A   i  �   i  �    �    �   i     i      �    �   i  c   i   	   D   !     �           '�       	   D   !     �       
�  '�  
�      _   ,      �      A  '�  A  '�  �      �      C  �    ����       U   �   U   �  �  Y  �  Y   U  �   U  �  5  �  5  �   U  ?   U  ?  5  �  5  �   U  
�   U  
�  5  1  5  1   U  �   U  �  5  y  5  y   U     U    5  �  5  �   U  _   U  _  5  	  5  	   U  �   U  �  5  Q  5  Q   U  �   U  �  5  �  5  �   U  7   U  7  5  �  5  �   U  !   U  !  5  ")  5  ")   U  $�   U  $�  5  %q  5  %q   U  '�   U  '�����    ����      C  �   �  �   �  
K      
K      
�  '�  
�  '�  
K  %q  
K  %q  +  $�  +  $�  
K  ")  
K  ")  +  !  +  !  
K  �  
K  �  +  7  +  7  
K  �  
K  �  +  �  +  �  
K  Q  
K  Q  +  �  +  �  
K  	  
K  	  +  _  +  _  
K  �  
K  �  +    +    
K  y  
K  y  +  �  +  �  
K  1  
K  1  +  
�  +  
�  
K  �  
K  �  +  ?  +  ?  
K  �  
K  �  +  �  +  �  
K  Y  
K  Y  �   �  �      C          �  
�  �  
�  �    �    	�  M  	�  M  O  K  O  K  	�  �  	�  �  O  �  O  �  	�  	�  	�  	�  O  1  O  1  �  $�  �  $�  3  1  3  1  �  	�  �  	�    �    �  �  �  �  �    K    K  �  M  �  M            C  �  �   �  �  �  %�  �  %�  �  �  �  �  	�  %  	�  %  O  #  O  #  	�  m  	�  m  O  k  O  k  	�  �  	�  �  O  �  O  �  	�  �  	�  �  O  �  O  �  	�  E  	�  E  O  C  O  C  	�  �  	�  �  O  �  O  �  	�   �  	�   �  O  "�  O  "�  	�  $  	�  $  O  &   O  &   	8  '3  	8  '3  m  &   m  &   �  $  �  $    "�    "�  �   �  �   �    �    �  �  �  �  �    C    C  �  E  �  E    �    �  �  �  �  �    �    �  �  �  �  �    e    e   �  �   �  �    k    k  �  m  �  m           �  s   �  s    #    #  �  %  �  %    �    �   �  �   �      C   ,   U  3   U  �  	�  �  	�  3   U  3      ^   ,      K      ^  '�  ^  '�  K      K      C  , ,   �  
K   �  
�  !�  
�  !�  
K   �  
K      C  , ,   �����   �   U  !�   U  !�����   �����      C  , ,   �  
K   �  
�  ;  
�  ;  
K   �  
K      C  , ,   �����   �   U  ;   U  ;����   �����      C  , ,  ]  
K  ]  
�    
�    
K  ]  
K      C  , ,  ]����  ]   U     U  ����  ]����      C  , ,  )  
K  )  
�  �  
�  �  
K  )  
K      C  , ,  )����  )   U  �   U  �����  )����      C  , ,  �  
K  �  
�  �  
�  �  
K  �  
K      C  , ,  �����  �   U  �   U  �����  �����      C  , ,  �  
K  �  
�  k  
�  k  
K  �  
K      C  , ,  �����  �   U  k   U  k����  �����      C  , ,  	�  
K  	�  
�  
7  
�  
7  
K  	�  
K      C  , ,  	�����  	�   U  
7   U  
7����  	�����      C  , ,  Y  
K  Y  
�    
�    
K  Y  
K      C  , ,  Y����  Y   U     U  ����  Y����      C  , ,  %  
K  %  
�  �  
�  �  
K  %  
K      C  , ,  %����  %   U  �   U  �����  %����      C  , ,  �  
K  �  
�  �  
�  �  
K  �  
K      C  , ,  �����  �   U  �   U  �����  �����      C  , ,  �  
K  �  
�  g  
�  g  
K  �  
K      C  , ,  �����  �   U  g   U  g����  �����      C  , ,  �  
K  �  
�  3  
�  3  
K  �  
K      C  , ,  �����  �   U  3   U  3����  �����      C  , ,  U  
K  U  
�  �  
�  �  
K  U  
K      C  , ,  U����  U   U  �   U  �����  U����      C  , ,  !  
K  !  
�  �  
�  �  
K  !  
K      C  , ,  !����  !   U  �   U  �����  !����      C  , ,  �  
K  �  
�  �  
�  �  
K  �  
K      C  , ,  �����  �   U  �   U  �����  �����      C  , ,  �  
K  �  
�  c  
�  c  
K  �  
K      C  , ,  �����  �   U  c   U  c����  �����      C  , ,  �  
K  �  
�  /  
�  /  
K  �  
K      C  , ,  �����  �   U  /   U  /����  �����      C  , ,  Q  
K  Q  
�  �  
�  �  
K  Q  
K      C  , ,  Q����  Q   U  �   U  �����  Q����      C  , ,    
K    
�  �  
�  �  
K    
K      C  , ,  ����     U  �   U  �����  ����      C  , ,  "�  
K  "�  
�  #_  
�  #_  
K  "�  
K      C  , ,  "�����  "�   U  #_   U  #_����  "�����      C  , ,  $�  
K  $�  
�  %+  
�  %+  
K  $�  
K      C  , ,  $�����  $�   U  %+   U  %+����  $�����      C  , ,  &M  
K  &M  
�  &�  
�  &�  
K  &M  
K      C  , ,  &M����  &M   U  &�   U  &�����  &M����      B  , ,  k  3  k  �    �    3  k  3      B  , ,  �  �  �  	[  e  	[  e  �  �  �      B  , ,  �  ]  �    e    e  ]  �  ]      B  , ,  �  	  �  �  e  �  e  	  �  	      B  , ,  �  �  �  9  e  9  e  �  �  �      B  , ,  �  ;  �  �  e  �  e  ;  �  ;      B  , ,  �  3  �  �  i  �  i  3  �  3      B  , ,  _  �  _  	y  	  	y  	  �  _  �      B  , ,  _  {  _  %  	  %  	  {  _  {      B  , ,  _  ;  _  �  	  �  	  ;  _  ;      B  , ,    3    �  �  �  �  3    3      B  , ,    �    	[  �  	[  �  �    �      B  , ,    ]      �    �  ]    ]      B  , ,    	    �  �  �  �  	    	      B  , ,    �    9  �  9  �  �    �      B  , ,    ;    �  �  �  �  ;    ;      B  , ,  g  3  g  �    �    3  g  3      B  , ,  �  �  �  	y  Q  	y  Q  �  �  �      B  , ,  �  {  �  %  Q  %  Q  {  �  {      B  , ,  �  ;  �  �  Q  �  Q  ;  �  ;      B  , ,  �  3  �  �  e  �  e  3  �  3      B  , ,    3    �  �  �  �  3    3      B  , ,  K  �  K  	[  �  	[  �  �  K  �      B  , ,  K  ]  K    �    �  ]  K  ]      B  , ,  K  	  K  �  �  �  �  	  K  	      B  , ,  K  �  K  9  �  9  �  �  K  �      B  , ,  K  ;  K  �  �  �  �  ;  K  ;      B  , ,  c  3  c  �    �    3  c  3      B  , ,  �  �  �  	y  �  	y  �  �  �  �      B  , ,  �  {  �  %  �  %  �  {  �  {      B  , ,  $�  ;  $�  �  %q  �  %q  ;  $�  ;      B  , ,  �  ;  �  �  �  �  �  ;  �  ;      B  , ,  �  3  �  �  a  �  a  3  �  3      B  , ,  �  �  �  	[  =  	[  =  �  �  �      B  , ,  �  ]  �    =    =  ]  �  ]      B  , ,  �  	  �  �  =  �  =  	  �  	      B  , ,  �  �  �  9  =  9  =  �  �  �      B  , ,  �  ;  �  �  =  �  =  ;  �  ;      B  , ,    3    �  �  �  �  3    3      B  , ,  7  �  7  	y  �  	y  �  �  7  �      B  , ,  7  {  7  %  �  %  �  {  7  {      B  , ,  7  ;  7  �  �  �  �  ;  7  ;      B  , ,  _  3  _  �  	  �  	  3  _  3      B  , ,  �  3  �  �   ]  �   ]  3  �  3      B  , ,  �  �  �  	[   �  	[   �  �  �  �      B  , ,  �  ]  �     �     �  ]  �  ]      B  , ,  �  	  �  �   �  �   �  	  �  	      B  , ,  �  �  �  9   �  9   �  �  �  �      B  , ,  �  ;  �  �   �  �   �  ;  �  ;      B  , ,  !  3  !  �  !�  �  !�  3  !  3      B  , ,  !  �  !  	y  ")  	y  ")  �  !  �      B  , ,  !  {  !  %  ")  %  ")  {  !  {      B  , ,  !  ;  !  �  ")  �  ")  ;  !  ;      B  , ,  "[  3  "[  �  #  �  #  3  "[  3      B  , ,  ##  �  ##  	[  #�  	[  #�  �  ##  �      B  , ,  ##  ]  ##    #�    #�  ]  ##  ]      B  , ,  ##  	  ##  �  #�  �  #�  	  ##  	      B  , ,  ##  �  ##  9  #�  9  #�  �  ##  �      B  , ,  ##  ;  ##  �  #�  �  #�  ;  ##  ;      B  , ,  #�  3  #�  �  $Y  �  $Y  3  #�  3      B  , ,  $�  �  $�  	y  %q  	y  %q  �  $�  �      B  , ,  $�  {  $�  %  %q  %  %q  {  $�  {      B  , ,  �  {  �  %  �  %  �  {  �  {      B  , ,  �  ;  �  �  �  �  �  ;  �  ;      B  , ,  �  3  �  �  U  �  U  3  �  3      B  , ,  �  �  �  	[  E  	[  E  �  �  �      B  , ,  ?  {  ?  %  �  %  �  {  ?  {      B  , ,  ?  ;  ?  �  �  �  �  ;  ?  ;      B  , ,  S  3  S  �  �  �  �  3  S  3      B  , ,  �  3  �  �  	Q  �  	Q  3  �  3      B  , ,  �  �  �  	[  	�  	[  	�  �  �  �      B  , ,  �  ]  �    	�    	�  ]  �  ]      B  , ,  �  	  �  �  	�  �  	�  	  �  	      B  , ,  �  �  �  9  	�  9  	�  �  �  �      B  , ,  �  ;  �  �  	�  �  	�  ;  �  ;      B  , ,  
�  �  
�  	y  1  	y  1  �  
�  �      B  , ,  s  ]  s          ]  s  ]      B  , ,  s  	  s  �    �    	  s  	      B  , ,  s  �  s  9    9    �  s  �      B  , ,  s  ;  s  �    �    ;  s  ;      B  , ,  �  3  �  �  m  �  m  3  �  3      B  , ,    �    	y  �  	y  �  �    �      B  , ,    {    %  �  %  �  {    {      B  , ,    3    �  �  �  �  3    3      B  , ,    ;    �  �  �  �  ;    ;      B  , ,  �  ]  �    E    E  ]  �  ]      B  , ,  �  	  �  �  E  �  E  	  �  	      B  , ,  �  �  �  9  E  9  E  �  �  �      B  , ,  �  ;  �  �  E  �  E  ;  �  ;      B  , ,  �  3  �  �  �  �  �  3  �  3      B  , ,  ?  �  ?  	y  �  	y  �  �  ?  �      B  , ,  S  ]  S    �    �  ]  S  ]      B  , ,  S  	  S  �  �  �  �  	  S  	      B  , ,  S  �  S  9  �  9  �  �  S  �      B  , ,  S  ;  S  �  �  �  �  ;  S  ;      B  , ,  W  3  W  �    �    3  W  3      B  , ,  �  �  �  	y  �  	y  �  �  �  �      B  , ,   �  �   �  	y  Y  	y  Y  �   �  �      B  , ,   �  {   �  %  Y  %  Y  {   �  {      B  , ,   �  '   �  �  Y  �  Y  '   �  '      B  , ,   �  �   �  9  Y  9  Y  �   �  �      B  , ,   �  ;   �  �  Y  �  Y  ;   �  ;      B  , ,    3    �  �  �  �  3    3      B  , ,  S  �  S  	[  �  	[  �  �  S  �      B  , ,  �  �  �  	y  y  	y  y  �  �  �      B  , ,  �  {  �  %  y  %  y  {  �  {      B  , ,  �  ;  �  �  y  �  y  ;  �  ;      B  , ,  o  3  o  �    �    3  o  3      B  , ,  s  �  s  	[    	[    �  s  �      B  , ,  
�  {  
�  %  1  %  1  {  
�  {      B  , ,  
�  ;  
�  �  1  �  1  ;  
�  ;      B  , ,  �  3  �  �  q  �  q  3  �  3      B  , ,  +  �  +  	[  �  	[  �  �  +  �      B  , ,  +  ]  +    �    �  ]  +  ]      B  , ,  +  	  +  �  �  �  �  	  +  	      B  , ,  +  �  +  9  �  9  �  �  +  �      B  , ,  +  ;  +  �  �  �  �  ;  +  ;      B  , ,    3    �  �  �  �  3    3      A   ,   �  �   �  	�  %�  	�  %�  �   �  �      A   ,   �   �   �  u  %�  u  %�   �   �   �      ]  , ,    ���B      �  '�  �  '����B    ���B      @   ,���B  ���B  ^  (F  ^  (F  ���B        D   ,   �����   �   U  @   U  @����   �����      D   ,   �  
K   �  
�  @  
�  @  
K   �  
K      �    ,              
�  '�  
�  '�                  z   ,   �����   �   U  @   U  @����   �����      @   ,   �  
K   �  
�  @  
�  @  
K   �  
K      C        @������     � A       C        @������   O  � A       C        @������   &�  � X       C        @������   &�  � X       @  ;      @������    �     VNB       @        @������    �  
� VPB       D        @������    �     VGND      D        @������    �  
� VPWR      Q   ,              
�  '�  
�  '�                  N  , ,      �      
�  '�  
�  '�  �      �      C   ,  �  Q  �  �  �  �  �  Q  �  Q      C   ,  �  Q  �  �  p  �  p  Q  �  Q      C   ,  &M  �  &M  O  &�  O  &�  �  &M  �      C   ,  &M  Q  &M  �  &�  �  &�  Q  &M  Q      S  ,    @������ BZ                
buf_16     � 
   % 0� 
   % 0 sky130_fd_sc_hd__buf_8    B   �  �   i  �  �   �  �   �    �    �  
7  !  
7  !    /    /  
7  �  
7  �    �    �  
7  i  
7  i   i  �   i  �    �    �   i  /   i  /    !    !   i  �   i      B  �  w   i  w  
7    
7            
7  �  
7  �    	�    	�  
7  
U  
7  
U    c    c  
7  �  
7  �          
7  �  
7  �    �    �  
7  A  
7  A    O    O  
7  �  
7  �    �    �  
7  �  
7  �   i  �   i  �    �    �   i  O   i  O    A    A   i  �   i  �    �    �   i     i      �    �   i  c   i  c    
U    
U   i  	�   i  	�    �    �   i     i             i  w   i   	   D   !     �       
�  �  
�   	   D   !     �           �          _   ,      �      A  �  A  �  �      �      C   �   �   �   �  �  �  �  �  �   _  �   _  	�  �  	�  �  O  �  O  �  	�  �  	�  �  O  ;  O  ;  �  �  �  �  3  ;  3  ;  �  �  �  �    �    �  �  Y  �  Y   �   �   �      C   �    ����       U     U    5  M  5  M   U  K   U  K  5  �  5  �   U  �   U  �  5  	�  5  	�   U  �   U  �  5  %  5  %   U  #   U  #  5  m  5  m   U  k   U  k  u  �  u  �   U  �   U  �����    ����      C   �  k  �  k  
K  m  
K  m  +  #  +  #  
K  %  
K  %  +  �  +  �  
K  	�  
K  	�  +  �  +  �  
K  E  
K  E  +  �  +  �  
K  �  
K  �  +  S  +  S  
K      
K      
�  �  
�  �  
K  �  
K  �  �  k  �      C    ?   �  ?  �  �  �  �  �  ?  �  ?  	�  �  	�  �  O  
�  O  
�  	�  1  	�  1  O  �  O  �  	�  y  	�  y  O    O    	�  �  	�  �   �     �    �  y  �  y   �  �   �  �  �  1  �  1   �  
�   �  
�  �  �  �  �   �  ?   �      C   ,   �  3   �  �  �  �  �  3   �  3      ^   ,      K      ^  �  ^  �  K      K      C  , ,   �  
K   �  
�  ;  
�  ;  
K   �  
K      C  , ,   �����   �   U  ;   U  ;����   �����      C  , ,  ]  
K  ]  
�    
�    
K  ]  
K      C  , ,  ]����  ]   U     U  ����  ]����      C  , ,  )  
K  )  
�  �  
�  �  
K  )  
K      C  , ,  )����  )   U  �   U  �����  )����      C  , ,  �  
K  �  
�  �  
�  �  
K  �  
K      C  , ,  �����  �   U  �   U  �����  �����      C  , ,  �  
K  �  
�  k  
�  k  
K  �  
K      C  , ,  �����  �   U  k   U  k����  �����      C  , ,  	�  
K  	�  
�  
7  
�  
7  
K  	�  
K      C  , ,  	�����  	�   U  
7   U  
7����  	�����      C  , ,  Y  
K  Y  
�    
�    
K  Y  
K      C  , ,  Y����  Y   U     U  ����  Y����      C  , ,  %  
K  %  
�  �  
�  �  
K  %  
K      C  , ,  %����  %   U  �   U  �����  %����      C  , ,  �  
K  �  
�  �  
�  �  
K  �  
K      C  , ,  �����  �   U  �   U  �����  �����      C  , ,  �  
K  �  
�  g  
�  g  
K  �  
K      C  , ,  �����  �   U  g   U  g����  �����      C  , ,  �  
K  �  
�  3  
�  3  
K  �  
K      C  , ,  �����  �   U  3   U  3����  �����      C  , ,  U  
K  U  
�  �  
�  �  
K  U  
K      C  , ,  U����  U   U  �   U  �����  U����      B  , ,  �  '  �  �  e  �  e  '  �  '      B  , ,  �  {  �  %  e  %  e  {  �  {      B  , ,  �  '  �  �  e  �  e  '  �  '      B  , ,  +  ;  +  �  �  �  �  ;  +  ;      B  , ,    3    �  )  �  )  3    3      B  , ,  �  �  �  0  y  0  y  �  �  �      B  , ,  �  �  �  �  y  �  y  �  �  �      B  , ,  +  {  +  %  �  %  �  {  +  {      B  , ,  
�  �  
�  0  1  0  1  �  
�  �      B  , ,  �  {  �  %  	�  %  	�  {  �  {      B  , ,  �  {  �  %  e  %  e  {  �  {      B  , ,  s  �  s  	y    	y    �  s  �      B  , ,  s  {  s  %    %    {  s  {      B  , ,  s  ;  s  �    �    ;  s  ;      B  , ,    a    	  �  	  �  a    a      B  , ,    �    0  �  0  �  �    �      B  , ,   �  �   �  	[  Y  	[  Y  �   �  �      B  , ,   �  ]   �    Y    Y  ]   �  ]      B  , ,   �  	   �  �  Y  �  Y  	   �  	      B  , ,   �  �   �  �  Y  �  Y  �   �  �      B  , ,   �  3   �  �  �  �  �  3   �  3      B  , ,  0  3  0  �  �  �  �  3  0  3      B  , ,  S  �  S  	y  �  	y  �  �  S  �      B  , ,  S  {  S  %  �  %  �  {  S  {      B  , ,  S  ;  S  �  �  �  �  ;  S  ;      B  , ,  �  3  �  �  .  �  .  3  �  3      B  , ,  �  �  �  	[  �  	[  �  �  �  �      B  , ,  �  ]  �    �    �  ]  �  ]      B  , ,  �  	  �  �  �  �  �  	  �  	      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  �  �  �  	y  E  	y  E  �  �  �      B  , ,  �  {  �  %  E  %  E  {  �  {      B  , ,  �  ;  �  �  E  �  E  ;  �  ;      B  , ,  �  3  �  �  �  �  �  3  �  3      B  , ,  ?  a  ?  	  �  	  �  a  ?  a      B  , ,  ?  �  ?  0  �  0  �  �  ?  �      B  , ,    �    �  �  �  �  �    �      B  , ,  �  �  �  	y  e  	y  e  �  �  �      B  , ,  ?  �  ?  �  �  �  �  �  ?  �      B  , ,  /  3  /  �  �  �  �  3  /  3      B  , ,  �  �  �  	y  	�  	y  	�  �  �  �      B  , ,  �  ;  �  �  	�  �  	�  ;  �  ;      B  , ,  	�  3  	�  �  
-  �  
-  3  	�  3      B  , ,  
�  a  
�  	  1  	  1  a  
�  a      B  , ,  
�  �  
�  �  1  �  1  �  
�  �      B  , ,  
�  3  
�  �  �  �  �  3  
�  3      B  , ,  +  �  +  	y  �  	y  �  �  +  �      B  , ,  +  3  +  �  �  �  �  3  +  3      B  , ,  �  3  �  �  }  �  }  3  �  3      B  , ,  �  a  �  	  y  	  y  a  �  a      A   ,   �  �   �  	�  �  	�  �  �   �  �      A   ,   �   �   �  u  �  u  �   �   �   �      ]  , ,    ���B      �  �  �  ����B    ���B      @   ,���B  ���B  ^  N  ^  N  ���B        D   ,   �����   �   U  @   U  @����   �����      D   ,   �  
K   �  
�  @  
�  @  
K   �  
K      �    ,              
�  �  
�  �                  z   ,   �����   �   U  @   U  @����   �����      @   ,   �  
K   �  
�  @  
�  @  
K   �  
K      C        @������   �  � A       C        @������     R X       C        @������     � X       C        @������   �  � A       C        @������    �     VGND      C        @������    �  
� VPWR      C        @������     � X       C        @������    �  � A       @  ;      @������    �     VNB       @        @������    �  
� VPB       D        @������    �     VGND      D        @������    �  
� VPWR      Q   ,              
�  �  
�  �                  N  , ,      �      
�  �  
�  �  �      �      C   ,   �  Q   �  �  @  �  @  Q   �  Q      C   ,  b  Q  b  �    �    Q  b  Q      C   ,  .  Q  .  �  �  �  �  Q  .  Q      C   ,  �  �  �  O  l  O  l  �  �  �      C   ,  �  Q  �  �  l  �  l  Q  �  Q      C   ,  �  �  �  �  l  �  l  �  �  �      C   ,   �����   �   U  @   U  @����   �����      C   ,   �  
K   �  
�  @  
�  @  
K   �  
K      S  ,    @������ BZ                
buf_8      � 
   % 0� 
   % 0 sky130_fd_sc_hd__buf_1    B   l  C   i  C  $  �  $  �  n  C  n  C  
7  �  
7  �  n  �  n  �  $  �  $  �   i  C   i      B   �  �   i  �  >  m  >  m  �   �  �   �  -  m  -  m  T  �  T  �  
7  !  
7  !  �    �    �  !  �  !   i  �   i   	   D   !     �           d       	   D   !     �       
�  d  
�      _   ,      �      �  d  �  d  �      �      C   L     �    �  [  �  [          	�    	�     �     �      C   L    ����       U     U    �  W  �  W   U  d   U  d����    ����      C   �   �   �   �  %  �  %  �  �   �  �   �  	�  Y  	�  Y  �  H  �  H  n  �  n  �  $  H  $  H  {  Y  {  Y   �   �   �      C   L    S    
K      
K      
�  d  
�  d  
K  W  
K  W  S    S      C   ,   i  �   i  K  �  K  �  �   i  �      ^   ,      �      ^  d  ^  d  �      �      C  , ,  )����  )   U  �   U  �����  )����      C  , ,  )  
K  )  
�  �  
�  �  
K  )  
K      C  , ,  ]����  ]   U     U  ����  ]����      C  , ,  ]  
K  ]  
�    
�    
K  ]  
K      C  , ,   �����   �   U  ;   U  ;����   �����      C  , ,   �  
K   �  
�  ;  
�  ;  
K   �  
K      B  , ,    �    g  �  g  �  �    �      B  , ,        �  �  �  �            B  , ,    �    	Q  �  	Q  �  �    �      B  , ,    t      �    �  t    t      B  , ,  ]  '  ]  �    �    '  ]  '      B  , ,  ]  S  ]  �    �    S  ]  S      B  , ,  ]  �  ]  	Q    	Q    �  ]  �      B  , ,   �  3   �  �  c  �  c  3   �  3      B  , ,   �  h   �    Y    Y  h   �  h      B  , ,   �  S   �  �  Y  �  Y  S   �  S      B  , ,   �  �   �  	Q  Y  	Q  Y  �   �  �      A   ,   �   �   �  �  �  �  �   �   �   �      A   ,   �  �   �  	�  �  	�  �  �   �  �      ]  , ,    ���B      �  d  �  d���B    ���B      @   ,���B  ���B  ^  "  ^  "  ���B        D   ,   �����   �   U  E   U  E����   �����      D   ,   �  
K   �  
�  ;  
�  ;  
K   �  
K      �    ,              
�  d  
�  d                  z   ,   �����   �   U  E   U  E����   �����      @   ,   �  
K   �  
�  ;  
�  ;  
K   �  
K      C        @������    �  
� VPWR      C        @������    �     VGND      C        @������   t  � X       C        @������   t  N X       C        @������   t  � X       C        @������    �  � A       @  ;      @������    �     VNB       @        @������    �  
� VPB       D        @������    �     VGND      D        @������    �  
� VPWR      Q   ,              
�  d  
�  d                  N  , ,      �      
�  d  
�  d  �      �      C   ,    �    S  �  S  �  �    �      C   ,    �    �  �  �  �  �    �      C   ,    M    �  �  �  �  M    M      C   ,   �  Q   �  �  ;  �  ;  Q   �  Q      C   ,   �  
K   �  
�  ;  
�  ;  
K   �  
K      C   ,   �����   �   U  E   U  E����   �����      S  ,    @������ BZ                
buf_1      � 
   % 0� 
   % 0 
pfet$6    B   ,  ����8  �  �  �  �  ����8  ����8      B   ,  �  �  �  �R  �  �R  �  �  �  �      A  , ,  �      �  �@  �  �@  �      �          D   ,   #   7   #  �	  �  �	  �   7   #   7      D   ,  �   7  �  �	  u  �	  u   7  �   7      D   ,  3  �:  3  �   e  �   e  �:  3  �:      _   ,  �  ��  �  �\  �  �\  �  ��  �  ��      C   ,   A   #   A  �  �  �  �   #   A   #      C   ,  �   #  �  �  W  �  W   #  �   #      C   ,    �X    �  y  �  y  �X    �X      C   ,  r   #  r  �  �  �  �   #  r   #      ^   ,������������  ��  �  ��  �������������      C  , ,   A  O3   A  O�   �  O�   �  O3   A  O3      C  , ,  �  O3  �  O�  S  O�  S  O3  �  O3      C  , ,    O3    O�  �  O�  �  O3    O3      C  , ,  �  O3  �  O�  �  O�  �  O3  �  O3      C  , ,  E  O3  E  O�  �  O�  �  O3  E  O3      C  , ,  �  O3  �  O�  W  O�  W  O3  �  O3      C  , ,   A  v�   A  w=   �  w=   �  v�   A  v�      C  , ,  �  v�  �  w=  S  w=  S  v�  �  v�      C  , ,    v�    w=  �  w=  �  v�    v�      C  , ,  �  v�  �  w=  �  w=  �  v�  �  v�      C  , ,  E  v�  E  w=  �  w=  �  v�  E  v�      C  , ,  �  v�  �  w=  W  w=  W  v�  �  v�      C  , ,  w  �X  w  �  !  �  !  �X  w  �X      C  , ,  �  |3  �  |�  �  |�  �  |3  �  |3      C  , ,  �  }�  �  ~E  �  ~E  �  }�  �  }�      C  , ,  �    �  �  �  �  �    �        C  , ,  �  �k  �  �  �  �  �  �k  �  �k      C  , ,  �  ��  �  �}  �  �}  �  ��  �  ��      C  , ,  �  �;  �  ��  �  ��  �  �;  �  �;      C  , ,  �  ��  �  �M  �  �M  �  ��  �  ��      C  , ,  �  �  �  ��  �  ��  �  �  �  �      C  , ,  �  �s  �  �  �  �  �  �s  �  �s      C  , ,  �  ��  �  ��  �  ��  �  ��  �  ��      C  , ,  �  �C  �  ��  �  ��  �  �C  �  �C      C  , ,  �  ��  �  �U  �  �U  �  ��  �  ��      C  , ,  �  �  �  ��  �  ��  �  �  �  �      C  , ,  �  �{  �  �%  �  �%  �  �{  �  �{      C  , ,  �  ��  �  ��  �  ��  �  ��  �  ��      C  , ,  �  �K  �  ��  �  ��  �  �K  �  �K      C  , ,  �  ��  �  �]  �  �]  �  ��  �  ��      C  , ,  �  �  �  ��  �  ��  �  �  �  �      C  , ,  �  ��  �  �-  �  �-  �  ��  �  ��      C  , ,  �  ��  �  ��  �  ��  �  ��  �  ��      C  , ,  �  �S  �  ��  �  ��  �  �S  �  �S      C  , ,  �  ��  �  �e  �  �e  �  ��  �  ��      C  , ,  �  �#  �  ��  �  ��  �  �#  �  �#      C  , ,  �  w�  �  x�  �  x�  �  w�  �  w�      C  , ,  E  w�  E  x�  �  x�  �  w�  E  w�      C  , ,  E  yc  E  z  �  z  �  yc  E  yc      C  , ,  E  z�  E  {u  �  {u  �  z�  E  z�      C  , ,  E  |3  E  |�  �  |�  �  |3  E  |3      C  , ,  E  }�  E  ~E  �  ~E  �  }�  E  }�      C  , ,  E    E  �  �  �  �    E        C  , ,  E  �k  E  �  �  �  �  �k  E  �k      C  , ,  E  ��  E  �}  �  �}  �  ��  E  ��      C  , ,  E  �;  E  ��  �  ��  �  �;  E  �;      C  , ,  E  ��  E  �M  �  �M  �  ��  E  ��      C  , ,  E  �  E  ��  �  ��  �  �  E  �      C  , ,  E  �s  E  �  �  �  �  �s  E  �s      C  , ,  E  ��  E  ��  �  ��  �  ��  E  ��      C  , ,  E  �C  E  ��  �  ��  �  �C  E  �C      C  , ,  E  ��  E  �U  �  �U  �  ��  E  ��      C  , ,  E  �  E  ��  �  ��  �  �  E  �      C  , ,  E  �{  E  �%  �  �%  �  �{  E  �{      C  , ,  E  ��  E  ��  �  ��  �  ��  E  ��      C  , ,  E  �K  E  ��  �  ��  �  �K  E  �K      C  , ,  E  ��  E  �]  �  �]  �  ��  E  ��      C  , ,  E  �  E  ��  �  ��  �  �  E  �      C  , ,  E  ��  E  �-  �  �-  �  ��  E  ��      C  , ,  E  ��  E  ��  �  ��  �  ��  E  ��      C  , ,  E  �S  E  ��  �  ��  �  �S  E  �S      C  , ,  E  ��  E  �e  �  �e  �  ��  E  ��      C  , ,  E  �#  E  ��  �  ��  �  �#  E  �#      C  , ,  �  yc  �  z  �  z  �  yc  �  yc      C  , ,  �  w�  �  x�  W  x�  W  w�  �  w�      C  , ,  �  yc  �  z  W  z  W  yc  �  yc      C  , ,  �  z�  �  {u  W  {u  W  z�  �  z�      C  , ,  �  |3  �  |�  W  |�  W  |3  �  |3      C  , ,  �  }�  �  ~E  W  ~E  W  }�  �  }�      C  , ,  �    �  �  W  �  W    �        C  , ,  �  �k  �  �  W  �  W  �k  �  �k      C  , ,  �  ��  �  �}  W  �}  W  ��  �  ��      C  , ,  �  �;  �  ��  W  ��  W  �;  �  �;      C  , ,  �  ��  �  �M  W  �M  W  ��  �  ��      C  , ,  �  �  �  ��  W  ��  W  �  �  �      C  , ,  �  �s  �  �  W  �  W  �s  �  �s      C  , ,  �  ��  �  ��  W  ��  W  ��  �  ��      C  , ,  �  �C  �  ��  W  ��  W  �C  �  �C      C  , ,  �  ��  �  �U  W  �U  W  ��  �  ��      C  , ,  �  �  �  ��  W  ��  W  �  �  �      C  , ,  �  �{  �  �%  W  �%  W  �{  �  �{      C  , ,  �  ��  �  ��  W  ��  W  ��  �  ��      C  , ,  �  �K  �  ��  W  ��  W  �K  �  �K      C  , ,  �  ��  �  �]  W  �]  W  ��  �  ��      C  , ,  �  �  �  ��  W  ��  W  �  �  �      C  , ,  �  ��  �  �-  W  �-  W  ��  �  ��      C  , ,  �  ��  �  ��  W  ��  W  ��  �  ��      C  , ,  �  �S  �  ��  W  ��  W  �S  �  �S      C  , ,  �  ��  �  �e  W  �e  W  ��  �  ��      C  , ,  �  �#  �  ��  W  ��  W  �#  �  �#      C  , ,  �  z�  �  {u  �  {u  �  z�  �  z�      C  , ,  �  �X  �  �  �  �  �  �X  �  �X      C  , ,  G  �X  G  �  �  �  �  �X  G  �X      C  , ,  �  �X  �  �  Y  �  Y  �X  �  �X      C  , ,    �X    �  �  �  �  �X    �X      C  , ,    �X    �  )  �  )  �X    �X      C  , ,   A  �s   A  �   �  �   �  �s   A  �s      C  , ,   A  ��   A  ��   �  ��   �  ��   A  ��      C  , ,   A  �C   A  ��   �  ��   �  �C   A  �C      C  , ,   A  ��   A  �U   �  �U   �  ��   A  ��      C  , ,   A  �   A  ��   �  ��   �  �   A  �      C  , ,   A  �{   A  �%   �  �%   �  �{   A  �{      C  , ,   A  ��   A  ��   �  ��   �  ��   A  ��      C  , ,   A  �K   A  ��   �  ��   �  �K   A  �K      C  , ,   A  ��   A  �]   �  �]   �  ��   A  ��      C  , ,   A  �   A  ��   �  ��   �  �   A  �      C  , ,   A  ��   A  �-   �  �-   �  ��   A  ��      C  , ,   A  ��   A  ��   �  ��   �  ��   A  ��      C  , ,   A  �S   A  ��   �  ��   �  �S   A  �S      C  , ,   A  ��   A  �e   �  �e   �  ��   A  ��      C  , ,   A  �#   A  ��   �  ��   �  �#   A  �#      C  , ,   A  w�   A  x�   �  x�   �  w�   A  w�      C  , ,  �  w�  �  x�  S  x�  S  w�  �  w�      C  , ,  �  yc  �  z  S  z  S  yc  �  yc      C  , ,  �  z�  �  {u  S  {u  S  z�  �  z�      C  , ,  �  |3  �  |�  S  |�  S  |3  �  |3      C  , ,  �  }�  �  ~E  S  ~E  S  }�  �  }�      C  , ,  �    �  �  S  �  S    �        C  , ,  �  �k  �  �  S  �  S  �k  �  �k      C  , ,  �  ��  �  �}  S  �}  S  ��  �  ��      C  , ,  �  �;  �  ��  S  ��  S  �;  �  �;      C  , ,  �  ��  �  �M  S  �M  S  ��  �  ��      C  , ,  �  �  �  ��  S  ��  S  �  �  �      C  , ,  �  �s  �  �  S  �  S  �s  �  �s      C  , ,  �  ��  �  ��  S  ��  S  ��  �  ��      C  , ,  �  �C  �  ��  S  ��  S  �C  �  �C      C  , ,  �  ��  �  �U  S  �U  S  ��  �  ��      C  , ,  �  �  �  ��  S  ��  S  �  �  �      C  , ,  �  �{  �  �%  S  �%  S  �{  �  �{      C  , ,  �  ��  �  ��  S  ��  S  ��  �  ��      C  , ,  �  �K  �  ��  S  ��  S  �K  �  �K      C  , ,  �  ��  �  �]  S  �]  S  ��  �  ��      C  , ,  �  �  �  ��  S  ��  S  �  �  �      C  , ,  �  ��  �  �-  S  �-  S  ��  �  ��      C  , ,  �  ��  �  ��  S  ��  S  ��  �  ��      C  , ,  �  �S  �  ��  S  ��  S  �S  �  �S      C  , ,  �  ��  �  �e  S  �e  S  ��  �  ��      C  , ,  �  �#  �  ��  S  ��  S  �#  �  �#      C  , ,   A  yc   A  z   �  z   �  yc   A  yc      C  , ,    w�    x�  �  x�  �  w�    w�      C  , ,    yc    z  �  z  �  yc    yc      C  , ,    z�    {u  �  {u  �  z�    z�      C  , ,    |3    |�  �  |�  �  |3    |3      C  , ,    }�    ~E  �  ~E  �  }�    }�      C  , ,        �  �  �  �            C  , ,    �k    �  �  �  �  �k    �k      C  , ,    ��    �}  �  �}  �  ��    ��      C  , ,    �;    ��  �  ��  �  �;    �;      C  , ,    ��    �M  �  �M  �  ��    ��      C  , ,    �    ��  �  ��  �  �    �      C  , ,    �s    �  �  �  �  �s    �s      C  , ,    ��    ��  �  ��  �  ��    ��      C  , ,    �C    ��  �  ��  �  �C    �C      C  , ,    ��    �U  �  �U  �  ��    ��      C  , ,    �    ��  �  ��  �  �    �      C  , ,    �{    �%  �  �%  �  �{    �{      C  , ,    ��    ��  �  ��  �  ��    ��      C  , ,    �K    ��  �  ��  �  �K    �K      C  , ,    ��    �]  �  �]  �  ��    ��      C  , ,    �    ��  �  ��  �  �    �      C  , ,    ��    �-  �  �-  �  ��    ��      C  , ,    ��    ��  �  ��  �  ��    ��      C  , ,    �S    ��  �  ��  �  �S    �S      C  , ,    ��    �e  �  �e  �  ��    ��      C  , ,    �#    ��  �  ��  �  �#    �#      C  , ,   A  z�   A  {u   �  {u   �  z�   A  z�      C  , ,   A  |3   A  |�   �  |�   �  |3   A  |3      C  , ,   A  }�   A  ~E   �  ~E   �  }�   A  }�      C  , ,  o  �X  o  �    �    �X  o  �X      C  , ,  �  �X  �  �  �  �  �  �X  �  �X      C  , ,  ?  �X  ?  �  �  �  �  �X  ?  �X      C  , ,  �  �X  �  �  	Q  �  	Q  �X  �  �X      C  , ,  
  �X  
  �  
�  �  
�  �X  
  �X      C  , ,   A     A  �   �  �   �     A        C  , ,   A  �k   A  �   �  �   �  �k   A  �k      C  , ,   A  ��   A  �}   �  �}   �  ��   A  ��      C  , ,   A  �;   A  ��   �  ��   �  �;   A  �;      C  , ,   A  ��   A  �M   �  �M   �  ��   A  ��      C  , ,   A  �   A  ��   �  ��   �  �   A  �      C  , ,   A  W�   A  XM   �  XM   �  W�   A  W�      C  , ,   A  Y   A  Y�   �  Y�   �  Y   A  Y      C  , ,   A  Zs   A  [   �  [   �  Zs   A  Zs      C  , ,   A  [�   A  \�   �  \�   �  [�   A  [�      C  , ,   A  ]C   A  ]�   �  ]�   �  ]C   A  ]C      C  , ,   A  P�   A  QE   �  QE   �  P�   A  P�      C  , ,  �  P�  �  QE  S  QE  S  P�  �  P�      C  , ,  �  R  �  R�  S  R�  S  R  �  R      C  , ,  �  Sk  �  T  S  T  S  Sk  �  Sk      C  , ,  �  T�  �  U}  S  U}  S  T�  �  T�      C  , ,   A  R   A  R�   �  R�   �  R   A  R      C  , ,    P�    QE  �  QE  �  P�    P�      C  , ,    R    R�  �  R�  �  R    R      C  , ,    Sk    T  �  T  �  Sk    Sk      C  , ,   A  T�   A  U}   �  U}   �  T�   A  T�      C  , ,    T�    U}  �  U}  �  T�    T�      C  , ,    V;    V�  �  V�  �  V;    V;      C  , ,    W�    XM  �  XM  �  W�    W�      C  , ,    Y    Y�  �  Y�  �  Y    Y      C  , ,    Zs    [  �  [  �  Zs    Zs      C  , ,    [�    \�  �  \�  �  [�    [�      C  , ,    ]C    ]�  �  ]�  �  ]C    ]C      C  , ,    ^�    _U  �  _U  �  ^�    ^�      C  , ,    `    `�  �  `�  �  `    `      C  , ,    a{    b%  �  b%  �  a{    a{      C  , ,    b�    c�  �  c�  �  b�    b�      C  , ,    dK    d�  �  d�  �  dK    dK      C  , ,    e�    f]  �  f]  �  e�    e�      C  , ,    g    g�  �  g�  �  g    g      C  , ,    h�    i-  �  i-  �  h�    h�      C  , ,    i�    j�  �  j�  �  i�    i�      C  , ,    kS    k�  �  k�  �  kS    kS      C  , ,    l�    me  �  me  �  l�    l�      C  , ,    n#    n�  �  n�  �  n#    n#      C  , ,    o�    p5  �  p5  �  o�    o�      C  , ,    p�    q�  �  q�  �  p�    p�      C  , ,    r[    s  �  s  �  r[    r[      C  , ,    s�    tm  �  tm  �  s�    s�      C  , ,    u+    u�  �  u�  �  u+    u+      C  , ,  �  V;  �  V�  S  V�  S  V;  �  V;      C  , ,  �  W�  �  XM  S  XM  S  W�  �  W�      C  , ,  �  Y  �  Y�  S  Y�  S  Y  �  Y      C  , ,   A  V;   A  V�   �  V�   �  V;   A  V;      C  , ,  �  Zs  �  [  S  [  S  Zs  �  Zs      C  , ,  �  [�  �  \�  S  \�  S  [�  �  [�      C  , ,  �  ]C  �  ]�  S  ]�  S  ]C  �  ]C      C  , ,  �  ^�  �  _U  S  _U  S  ^�  �  ^�      C  , ,  �  `  �  `�  S  `�  S  `  �  `      C  , ,  �  a{  �  b%  S  b%  S  a{  �  a{      C  , ,  �  b�  �  c�  S  c�  S  b�  �  b�      C  , ,  �  dK  �  d�  S  d�  S  dK  �  dK      C  , ,  �  e�  �  f]  S  f]  S  e�  �  e�      C  , ,  �  g  �  g�  S  g�  S  g  �  g      C  , ,  �  h�  �  i-  S  i-  S  h�  �  h�      C  , ,  �  i�  �  j�  S  j�  S  i�  �  i�      C  , ,  �  kS  �  k�  S  k�  S  kS  �  kS      C  , ,  �  l�  �  me  S  me  S  l�  �  l�      C  , ,  �  n#  �  n�  S  n�  S  n#  �  n#      C  , ,  �  o�  �  p5  S  p5  S  o�  �  o�      C  , ,  �  p�  �  q�  S  q�  S  p�  �  p�      C  , ,  �  r[  �  s  S  s  S  r[  �  r[      C  , ,  �  s�  �  tm  S  tm  S  s�  �  s�      C  , ,  �  u+  �  u�  S  u�  S  u+  �  u+      C  , ,   A  ^�   A  _U   �  _U   �  ^�   A  ^�      C  , ,   A  `   A  `�   �  `�   �  `   A  `      C  , ,   A  a{   A  b%   �  b%   �  a{   A  a{      C  , ,   A  b�   A  c�   �  c�   �  b�   A  b�      C  , ,   A  Sk   A  T   �  T   �  Sk   A  Sk      C  , ,   A  dK   A  d�   �  d�   �  dK   A  dK      C  , ,   A  e�   A  f]   �  f]   �  e�   A  e�      C  , ,   A  g   A  g�   �  g�   �  g   A  g      C  , ,   A  h�   A  i-   �  i-   �  h�   A  h�      C  , ,   A  i�   A  j�   �  j�   �  i�   A  i�      C  , ,   A  kS   A  k�   �  k�   �  kS   A  kS      C  , ,   A  l�   A  me   �  me   �  l�   A  l�      C  , ,   A  n#   A  n�   �  n�   �  n#   A  n#      C  , ,   A  o�   A  p5   �  p5   �  o�   A  o�      C  , ,   A  p�   A  q�   �  q�   �  p�   A  p�      C  , ,   A  r[   A  s   �  s   �  r[   A  r[      C  , ,   A  s�   A  tm   �  tm   �  s�   A  s�      C  , ,   A  u+   A  u�   �  u�   �  u+   A  u+      C  , ,  �  b�  �  c�  �  c�  �  b�  �  b�      C  , ,  �  dK  �  d�  �  d�  �  dK  �  dK      C  , ,  �  e�  �  f]  �  f]  �  e�  �  e�      C  , ,  �  g  �  g�  �  g�  �  g  �  g      C  , ,  �  h�  �  i-  �  i-  �  h�  �  h�      C  , ,  �  i�  �  j�  �  j�  �  i�  �  i�      C  , ,  �  kS  �  k�  �  k�  �  kS  �  kS      C  , ,  �  l�  �  me  �  me  �  l�  �  l�      C  , ,  �  n#  �  n�  �  n�  �  n#  �  n#      C  , ,  �  o�  �  p5  �  p5  �  o�  �  o�      C  , ,  �  p�  �  q�  �  q�  �  p�  �  p�      C  , ,  �  r[  �  s  �  s  �  r[  �  r[      C  , ,  �  s�  �  tm  �  tm  �  s�  �  s�      C  , ,  �  u+  �  u�  �  u�  �  u+  �  u+      C  , ,  �  P�  �  QE  �  QE  �  P�  �  P�      C  , ,  E  P�  E  QE  �  QE  �  P�  E  P�      C  , ,  �  P�  �  QE  W  QE  W  P�  �  P�      C  , ,  �  R  �  R�  W  R�  W  R  �  R      C  , ,  �  Sk  �  T  W  T  W  Sk  �  Sk      C  , ,  �  T�  �  U}  W  U}  W  T�  �  T�      C  , ,  �  V;  �  V�  W  V�  W  V;  �  V;      C  , ,  �  W�  �  XM  W  XM  W  W�  �  W�      C  , ,  �  Y  �  Y�  W  Y�  W  Y  �  Y      C  , ,  �  Zs  �  [  W  [  W  Zs  �  Zs      C  , ,  �  [�  �  \�  W  \�  W  [�  �  [�      C  , ,  �  ]C  �  ]�  W  ]�  W  ]C  �  ]C      C  , ,  �  ^�  �  _U  W  _U  W  ^�  �  ^�      C  , ,  �  `  �  `�  W  `�  W  `  �  `      C  , ,  �  a{  �  b%  W  b%  W  a{  �  a{      C  , ,  �  b�  �  c�  W  c�  W  b�  �  b�      C  , ,  �  dK  �  d�  W  d�  W  dK  �  dK      C  , ,  �  e�  �  f]  W  f]  W  e�  �  e�      C  , ,  �  g  �  g�  W  g�  W  g  �  g      C  , ,  �  h�  �  i-  W  i-  W  h�  �  h�      C  , ,  �  i�  �  j�  W  j�  W  i�  �  i�      C  , ,  �  kS  �  k�  W  k�  W  kS  �  kS      C  , ,  �  l�  �  me  W  me  W  l�  �  l�      C  , ,  �  n#  �  n�  W  n�  W  n#  �  n#      C  , ,  �  o�  �  p5  W  p5  W  o�  �  o�      C  , ,  �  p�  �  q�  W  q�  W  p�  �  p�      C  , ,  �  r[  �  s  W  s  W  r[  �  r[      C  , ,  �  s�  �  tm  W  tm  W  s�  �  s�      C  , ,  �  u+  �  u�  W  u�  W  u+  �  u+      C  , ,  E  R  E  R�  �  R�  �  R  E  R      C  , ,  E  Sk  E  T  �  T  �  Sk  E  Sk      C  , ,  E  T�  E  U}  �  U}  �  T�  E  T�      C  , ,  E  V;  E  V�  �  V�  �  V;  E  V;      C  , ,  E  W�  E  XM  �  XM  �  W�  E  W�      C  , ,  E  Y  E  Y�  �  Y�  �  Y  E  Y      C  , ,  E  Zs  E  [  �  [  �  Zs  E  Zs      C  , ,  E  [�  E  \�  �  \�  �  [�  E  [�      C  , ,  E  ]C  E  ]�  �  ]�  �  ]C  E  ]C      C  , ,  E  ^�  E  _U  �  _U  �  ^�  E  ^�      C  , ,  E  `  E  `�  �  `�  �  `  E  `      C  , ,  E  a{  E  b%  �  b%  �  a{  E  a{      C  , ,  E  b�  E  c�  �  c�  �  b�  E  b�      C  , ,  E  dK  E  d�  �  d�  �  dK  E  dK      C  , ,  E  e�  E  f]  �  f]  �  e�  E  e�      C  , ,  E  g  E  g�  �  g�  �  g  E  g      C  , ,  E  h�  E  i-  �  i-  �  h�  E  h�      C  , ,  E  i�  E  j�  �  j�  �  i�  E  i�      C  , ,  E  kS  E  k�  �  k�  �  kS  E  kS      C  , ,  E  l�  E  me  �  me  �  l�  E  l�      C  , ,  E  n#  E  n�  �  n�  �  n#  E  n#      C  , ,  E  o�  E  p5  �  p5  �  o�  E  o�      C  , ,  E  p�  E  q�  �  q�  �  p�  E  p�      C  , ,  E  r[  E  s  �  s  �  r[  E  r[      C  , ,  E  s�  E  tm  �  tm  �  s�  E  s�      C  , ,  E  u+  E  u�  �  u�  �  u+  E  u+      C  , ,  �  R  �  R�  �  R�  �  R  �  R      C  , ,  �  Sk  �  T  �  T  �  Sk  �  Sk      C  , ,  �  T�  �  U}  �  U}  �  T�  �  T�      C  , ,  �  V;  �  V�  �  V�  �  V;  �  V;      C  , ,  �  W�  �  XM  �  XM  �  W�  �  W�      C  , ,  �  Y  �  Y�  �  Y�  �  Y  �  Y      C  , ,  �  Zs  �  [  �  [  �  Zs  �  Zs      C  , ,  �  [�  �  \�  �  \�  �  [�  �  [�      C  , ,  �  ]C  �  ]�  �  ]�  �  ]C  �  ]C      C  , ,  �  ^�  �  _U  �  _U  �  ^�  �  ^�      C  , ,  �  `  �  `�  �  `�  �  `  �  `      C  , ,  �  a{  �  b%  �  b%  �  a{  �  a{      C  , ,  �  '�  �  (}  �  (}  �  '�  �  '�      C  , ,   A  '�   A  (}   �  (}   �  '�   A  '�      C  , ,  E  '�  E  (}  �  (}  �  '�  E  '�      C  , ,    '�    (}  �  (}  �  '�    '�      C  , ,  �  '�  �  (}  W  (}  W  '�  �  '�      C  , ,  �  '�  �  (}  S  (}  S  '�  �  '�      C  , ,  �  0C  �  0�  �  0�  �  0C  �  0C      C  , ,  �  1�  �  2U  �  2U  �  1�  �  1�      C  , ,  �  3  �  3�  �  3�  �  3  �  3      C  , ,  �  4{  �  5%  �  5%  �  4{  �  4{      C  , ,  �  5�  �  6�  �  6�  �  5�  �  5�      C  , ,  �  7K  �  7�  �  7�  �  7K  �  7K      C  , ,  �  8�  �  9]  �  9]  �  8�  �  8�      C  , ,  �  :  �  :�  �  :�  �  :  �  :      C  , ,  �  ;�  �  <-  �  <-  �  ;�  �  ;�      C  , ,  �  <�  �  =�  �  =�  �  <�  �  <�      C  , ,  �  >S  �  >�  �  >�  �  >S  �  >S      C  , ,  �  ?�  �  @e  �  @e  �  ?�  �  ?�      C  , ,  �  A#  �  A�  �  A�  �  A#  �  A#      C  , ,  �  B�  �  C5  �  C5  �  B�  �  B�      C  , ,  �  C�  �  D�  �  D�  �  C�  �  C�      C  , ,  �  E[  �  F  �  F  �  E[  �  E[      C  , ,  �  F�  �  Gm  �  Gm  �  F�  �  F�      C  , ,  �  H+  �  H�  �  H�  �  H+  �  H+      C  , ,  �  I�  �  J=  �  J=  �  I�  �  I�      C  , ,  �  J�  �  K�  �  K�  �  J�  �  J�      C  , ,  �  Lc  �  M  �  M  �  Lc  �  Lc      C  , ,  �  M�  �  Nu  �  Nu  �  M�  �  M�      C  , ,  �  );  �  )�  �  )�  �  );  �  );      C  , ,  �  *�  �  +M  �  +M  �  *�  �  *�      C  , ,  E  );  E  )�  �  )�  �  );  E  );      C  , ,  E  *�  E  +M  �  +M  �  *�  E  *�      C  , ,  E  ,  E  ,�  �  ,�  �  ,  E  ,      C  , ,  E  -s  E  .  �  .  �  -s  E  -s      C  , ,  E  .�  E  /�  �  /�  �  .�  E  .�      C  , ,  E  0C  E  0�  �  0�  �  0C  E  0C      C  , ,  E  1�  E  2U  �  2U  �  1�  E  1�      C  , ,  E  3  E  3�  �  3�  �  3  E  3      C  , ,  E  4{  E  5%  �  5%  �  4{  E  4{      C  , ,  E  5�  E  6�  �  6�  �  5�  E  5�      C  , ,  E  7K  E  7�  �  7�  �  7K  E  7K      C  , ,  E  8�  E  9]  �  9]  �  8�  E  8�      C  , ,  E  :  E  :�  �  :�  �  :  E  :      C  , ,  E  ;�  E  <-  �  <-  �  ;�  E  ;�      C  , ,  E  <�  E  =�  �  =�  �  <�  E  <�      C  , ,  E  >S  E  >�  �  >�  �  >S  E  >S      C  , ,  E  ?�  E  @e  �  @e  �  ?�  E  ?�      C  , ,  E  A#  E  A�  �  A�  �  A#  E  A#      C  , ,  E  B�  E  C5  �  C5  �  B�  E  B�      C  , ,  E  C�  E  D�  �  D�  �  C�  E  C�      C  , ,  E  E[  E  F  �  F  �  E[  E  E[      C  , ,  E  F�  E  Gm  �  Gm  �  F�  E  F�      C  , ,  E  H+  E  H�  �  H�  �  H+  E  H+      C  , ,  E  I�  E  J=  �  J=  �  I�  E  I�      C  , ,  E  J�  E  K�  �  K�  �  J�  E  J�      C  , ,  E  Lc  E  M  �  M  �  Lc  E  Lc      C  , ,  E  M�  E  Nu  �  Nu  �  M�  E  M�      C  , ,  �  ,  �  ,�  �  ,�  �  ,  �  ,      C  , ,  �  -s  �  .  �  .  �  -s  �  -s      C  , ,  �  );  �  )�  W  )�  W  );  �  );      C  , ,  �  *�  �  +M  W  +M  W  *�  �  *�      C  , ,  �  ,  �  ,�  W  ,�  W  ,  �  ,      C  , ,  �  -s  �  .  W  .  W  -s  �  -s      C  , ,  �  .�  �  /�  W  /�  W  .�  �  .�      C  , ,  �  0C  �  0�  W  0�  W  0C  �  0C      C  , ,  �  1�  �  2U  W  2U  W  1�  �  1�      C  , ,  �  3  �  3�  W  3�  W  3  �  3      C  , ,  �  4{  �  5%  W  5%  W  4{  �  4{      C  , ,  �  5�  �  6�  W  6�  W  5�  �  5�      C  , ,  �  7K  �  7�  W  7�  W  7K  �  7K      C  , ,  �  8�  �  9]  W  9]  W  8�  �  8�      C  , ,  �  :  �  :�  W  :�  W  :  �  :      C  , ,  �  ;�  �  <-  W  <-  W  ;�  �  ;�      C  , ,  �  <�  �  =�  W  =�  W  <�  �  <�      C  , ,  �  >S  �  >�  W  >�  W  >S  �  >S      C  , ,  �  ?�  �  @e  W  @e  W  ?�  �  ?�      C  , ,  �  A#  �  A�  W  A�  W  A#  �  A#      C  , ,  �  B�  �  C5  W  C5  W  B�  �  B�      C  , ,  �  C�  �  D�  W  D�  W  C�  �  C�      C  , ,  �  E[  �  F  W  F  W  E[  �  E[      C  , ,  �  F�  �  Gm  W  Gm  W  F�  �  F�      C  , ,  �  H+  �  H�  W  H�  W  H+  �  H+      C  , ,  �  I�  �  J=  W  J=  W  I�  �  I�      C  , ,  �  J�  �  K�  W  K�  W  J�  �  J�      C  , ,  �  Lc  �  M  W  M  W  Lc  �  Lc      C  , ,  �  M�  �  Nu  W  Nu  W  M�  �  M�      C  , ,  �  .�  �  /�  �  /�  �  .�  �  .�      C  , ,    *�    +M  �  +M  �  *�    *�      C  , ,    ,    ,�  �  ,�  �  ,    ,      C  , ,    -s    .  �  .  �  -s    -s      C  , ,    .�    /�  �  /�  �  .�    .�      C  , ,    0C    0�  �  0�  �  0C    0C      C  , ,    1�    2U  �  2U  �  1�    1�      C  , ,    3    3�  �  3�  �  3    3      C  , ,    4{    5%  �  5%  �  4{    4{      C  , ,    5�    6�  �  6�  �  5�    5�      C  , ,    7K    7�  �  7�  �  7K    7K      C  , ,    8�    9]  �  9]  �  8�    8�      C  , ,    :    :�  �  :�  �  :    :      C  , ,    ;�    <-  �  <-  �  ;�    ;�      C  , ,    <�    =�  �  =�  �  <�    <�      C  , ,    >S    >�  �  >�  �  >S    >S      C  , ,    ?�    @e  �  @e  �  ?�    ?�      C  , ,    A#    A�  �  A�  �  A#    A#      C  , ,    B�    C5  �  C5  �  B�    B�      C  , ,    C�    D�  �  D�  �  C�    C�      C  , ,    E[    F  �  F  �  E[    E[      C  , ,    F�    Gm  �  Gm  �  F�    F�      C  , ,    H+    H�  �  H�  �  H+    H+      C  , ,    I�    J=  �  J=  �  I�    I�      C  , ,   A  );   A  )�   �  )�   �  );   A  );      C  , ,   A  *�   A  +M   �  +M   �  *�   A  *�      C  , ,   A  ,   A  ,�   �  ,�   �  ,   A  ,      C  , ,   A  -s   A  .   �  .   �  -s   A  -s      C  , ,   A  .�   A  /�   �  /�   �  .�   A  .�      C  , ,   A  0C   A  0�   �  0�   �  0C   A  0C      C  , ,   A  1�   A  2U   �  2U   �  1�   A  1�      C  , ,   A  3   A  3�   �  3�   �  3   A  3      C  , ,   A  4{   A  5%   �  5%   �  4{   A  4{      C  , ,   A  5�   A  6�   �  6�   �  5�   A  5�      C  , ,   A  7K   A  7�   �  7�   �  7K   A  7K      C  , ,   A  8�   A  9]   �  9]   �  8�   A  8�      C  , ,   A  :   A  :�   �  :�   �  :   A  :      C  , ,   A  ;�   A  <-   �  <-   �  ;�   A  ;�      C  , ,   A  <�   A  =�   �  =�   �  <�   A  <�      C  , ,   A  >S   A  >�   �  >�   �  >S   A  >S      C  , ,   A  ?�   A  @e   �  @e   �  ?�   A  ?�      C  , ,   A  A#   A  A�   �  A�   �  A#   A  A#      C  , ,   A  B�   A  C5   �  C5   �  B�   A  B�      C  , ,   A  C�   A  D�   �  D�   �  C�   A  C�      C  , ,   A  E[   A  F   �  F   �  E[   A  E[      C  , ,   A  F�   A  Gm   �  Gm   �  F�   A  F�      C  , ,   A  H+   A  H�   �  H�   �  H+   A  H+      C  , ,  �  M�  �  Nu  S  Nu  S  M�  �  M�      C  , ,   A  M�   A  Nu   �  Nu   �  M�   A  M�      C  , ,   A  I�   A  J=   �  J=   �  I�   A  I�      C  , ,   A  J�   A  K�   �  K�   �  J�   A  J�      C  , ,  �  Lc  �  M  S  M  S  Lc  �  Lc      C  , ,    J�    K�  �  K�  �  J�    J�      C  , ,    Lc    M  �  M  �  Lc    Lc      C  , ,    M�    Nu  �  Nu  �  M�    M�      C  , ,   A  Lc   A  M   �  M   �  Lc   A  Lc      C  , ,    );    )�  �  )�  �  );    );      C  , ,  �  );  �  )�  S  )�  S  );  �  );      C  , ,  �  *�  �  +M  S  +M  S  *�  �  *�      C  , ,  �  ,  �  ,�  S  ,�  S  ,  �  ,      C  , ,  �  -s  �  .  S  .  S  -s  �  -s      C  , ,  �  .�  �  /�  S  /�  S  .�  �  .�      C  , ,  �  0C  �  0�  S  0�  S  0C  �  0C      C  , ,  �  1�  �  2U  S  2U  S  1�  �  1�      C  , ,  �  3  �  3�  S  3�  S  3  �  3      C  , ,  �  4{  �  5%  S  5%  S  4{  �  4{      C  , ,  �  5�  �  6�  S  6�  S  5�  �  5�      C  , ,  �  7K  �  7�  S  7�  S  7K  �  7K      C  , ,  �  8�  �  9]  S  9]  S  8�  �  8�      C  , ,  �  :  �  :�  S  :�  S  :  �  :      C  , ,  �  ;�  �  <-  S  <-  S  ;�  �  ;�      C  , ,  �  <�  �  =�  S  =�  S  <�  �  <�      C  , ,  �  >S  �  >�  S  >�  S  >S  �  >S      C  , ,  �  ?�  �  @e  S  @e  S  ?�  �  ?�      C  , ,  �  A#  �  A�  S  A�  S  A#  �  A#      C  , ,  �  B�  �  C5  S  C5  S  B�  �  B�      C  , ,  �  C�  �  D�  S  D�  S  C�  �  C�      C  , ,  �  E[  �  F  S  F  S  E[  �  E[      C  , ,  �  F�  �  Gm  S  Gm  S  F�  �  F�      C  , ,  �  H+  �  H�  S  H�  S  H+  �  H+      C  , ,  �  I�  �  J=  S  J=  S  I�  �  I�      C  , ,  �  J�  �  K�  S  K�  S  J�  �  J�      C  , ,   A  #�   A  $E   �  $E   �  #�   A  #�      C  , ,     s      �    �   s     s      C  , ,    �    �  �  �  �  �    �      C  , ,    C    �  �  �  �  C    C      C  , ,    �    U  �  U  �  �    �      C  , ,        �  �  �  �            C  , ,    {    %  �  %  �  {    {      C  , ,    �    	�  �  	�  �  �    �      C  , ,    
K    
�  �  
�  �  
K    
K      C  , ,    �    ]  �  ]  �  �    �      C  , ,        �  �  �  �            C  , ,    �    -  �  -  �  �    �      C  , ,    �    �  �  �  �  �    �      C  , ,    S    �  �  �  �  S    S      C  , ,    �    e  �  e  �  �    �      C  , ,    #    �  �  �  �  #    #      C  , ,    �    5  �  5  �  �    �      C  , ,    �    �  �  �  �  �    �      C  , ,    [      �    �  [    [      C  , ,    �    m  �  m  �  �    �      C  , ,    +    �  �  �  �  +    +      C  , ,    �    =  �  =  �  �    �      C  , ,    �    �  �  �  �  �    �      C  , ,    c       �     �  c    c      C  , ,     �    !u  �  !u  �   �     �      C  , ,    "3    "�  �  "�  �  "3    "3      C  , ,    #�    $E  �  $E  �  #�    #�      C  , ,    %    %�  �  %�  �  %    %      C  , ,    &k    '  �  '  �  &k    &k      C  , ,   A  %   A  %�   �  %�   �  %   A  %      C  , ,  �   s  �    S    S   s  �   s      C  , ,  �  �  �  �  S  �  S  �  �  �      C  , ,  �  C  �  �  S  �  S  C  �  C      C  , ,  �  �  �  U  S  U  S  �  �  �      C  , ,  �    �  �  S  �  S    �        C  , ,  �  {  �  %  S  %  S  {  �  {      C  , ,  �  �  �  	�  S  	�  S  �  �  �      C  , ,  �  
K  �  
�  S  
�  S  
K  �  
K      C  , ,  �  �  �  ]  S  ]  S  �  �  �      C  , ,  �    �  �  S  �  S    �        C  , ,  �  �  �  -  S  -  S  �  �  �      C  , ,  �  �  �  �  S  �  S  �  �  �      C  , ,  �  S  �  �  S  �  S  S  �  S      C  , ,  �  �  �  e  S  e  S  �  �  �      C  , ,  �  #  �  �  S  �  S  #  �  #      C  , ,  �  �  �  5  S  5  S  �  �  �      C  , ,  �  �  �  �  S  �  S  �  �  �      C  , ,  �  [  �    S    S  [  �  [      C  , ,  �  �  �  m  S  m  S  �  �  �      C  , ,  �  +  �  �  S  �  S  +  �  +      C  , ,  �  �  �  =  S  =  S  �  �  �      C  , ,  �  �  �  �  S  �  S  �  �  �      C  , ,  �  c  �     S     S  c  �  c      C  , ,  �   �  �  !u  S  !u  S   �  �   �      C  , ,  �  "3  �  "�  S  "�  S  "3  �  "3      C  , ,  �  #�  �  $E  S  $E  S  #�  �  #�      C  , ,  �  %  �  %�  S  %�  S  %  �  %      C  , ,  �  &k  �  '  S  '  S  &k  �  &k      C  , ,   A  &k   A  '   �  '   �  &k   A  &k      C  , ,   A   s   A     �     �   s   A   s      C  , ,   A  �   A  �   �  �   �  �   A  �      C  , ,   A  C   A  �   �  �   �  C   A  C      C  , ,   A  �   A  U   �  U   �  �   A  �      C  , ,   A     A  �   �  �   �     A        C  , ,   A  {   A  %   �  %   �  {   A  {      C  , ,   A  �   A  	�   �  	�   �  �   A  �      C  , ,   A  
K   A  
�   �  
�   �  
K   A  
K      C  , ,   A  �   A  ]   �  ]   �  �   A  �      C  , ,   A     A  �   �  �   �     A        C  , ,   A  �   A  -   �  -   �  �   A  �      C  , ,   A  �   A  �   �  �   �  �   A  �      C  , ,   A  S   A  �   �  �   �  S   A  S      C  , ,   A  �   A  e   �  e   �  �   A  �      C  , ,   A  #   A  �   �  �   �  #   A  #      C  , ,   A  �   A  5   �  5   �  �   A  �      C  , ,   A  �   A  �   �  �   �  �   A  �      C  , ,   A  [   A     �     �  [   A  [      C  , ,   A  �   A  m   �  m   �  �   A  �      C  , ,   A  +   A  �   �  �   �  +   A  +      C  , ,   A  �   A  =   �  =   �  �   A  �      C  , ,   A  �   A  �   �  �   �  �   A  �      C  , ,   A  c   A      �      �  c   A  c      C  , ,   A   �   A  !u   �  !u   �   �   A   �      C  , ,   A  "3   A  "�   �  "�   �  "3   A  "3      C  , ,  E  #�  E  $E  �  $E  �  #�  E  #�      C  , ,  E  %  E  %�  �  %�  �  %  E  %      C  , ,  E  &k  E  '  �  '  �  &k  E  &k      C  , ,  �  �  �  �  �  �  �  �  �  �      C  , ,  �  S  �  �  �  �  �  S  �  S      C  , ,  �  �  �  e  �  e  �  �  �  �      C  , ,  �  #  �  �  �  �  �  #  �  #      C  , ,  �  �  �  5  �  5  �  �  �  �      C  , ,  �  �  �  �  �  �  �  �  �  �      C  , ,  �  [  �    �    �  [  �  [      C  , ,  �  �  �  m  �  m  �  �  �  �      C  , ,  �  +  �  �  �  �  �  +  �  +      C  , ,  �  �  �  =  �  =  �  �  �  �      C  , ,  �  �  �  �  �  �  �  �  �  �      C  , ,  �  c  �     �     �  c  �  c      C  , ,  �   �  �  !u  �  !u  �   �  �   �      C  , ,  �  "3  �  "�  �  "�  �  "3  �  "3      C  , ,  �  #�  �  $E  �  $E  �  #�  �  #�      C  , ,  �  %  �  %�  �  %�  �  %  �  %      C  , ,  �  &k  �  '  �  '  �  &k  �  &k      C  , ,  �  �  �  ]  �  ]  �  �  �  �      C  , ,  �    �  �  �  �  �    �        C  , ,  �  �  �  -  �  -  �  �  �  �      C  , ,  E   s  E    �    �   s  E   s      C  , ,  E  �  E  �  �  �  �  �  E  �      C  , ,  E  C  E  �  �  �  �  C  E  C      C  , ,  E  �  E  U  �  U  �  �  E  �      C  , ,  E    E  �  �  �  �    E        C  , ,  E  {  E  %  �  %  �  {  E  {      C  , ,  E  �  E  	�  �  	�  �  �  E  �      C  , ,  E  
K  E  
�  �  
�  �  
K  E  
K      C  , ,  E  �  E  ]  �  ]  �  �  E  �      C  , ,  E    E  �  �  �  �    E        C  , ,  E  �  E  -  �  -  �  �  E  �      C  , ,  E  �  E  �  �  �  �  �  E  �      C  , ,  E  S  E  �  �  �  �  S  E  S      C  , ,  E  �  E  e  �  e  �  �  E  �      C  , ,  E  #  E  �  �  �  �  #  E  #      C  , ,  �   s  �    W    W   s  �   s      C  , ,  �  �  �  �  W  �  W  �  �  �      C  , ,  �  C  �  �  W  �  W  C  �  C      C  , ,  �  �  �  U  W  U  W  �  �  �      C  , ,  �    �  �  W  �  W    �        C  , ,  �  {  �  %  W  %  W  {  �  {      C  , ,  �  �  �  	�  W  	�  W  �  �  �      C  , ,  �  
K  �  
�  W  
�  W  
K  �  
K      C  , ,  �  �  �  ]  W  ]  W  �  �  �      C  , ,  �    �  �  W  �  W    �        C  , ,  �  �  �  -  W  -  W  �  �  �      C  , ,  �  �  �  �  W  �  W  �  �  �      C  , ,  �  S  �  �  W  �  W  S  �  S      C  , ,  �  �  �  e  W  e  W  �  �  �      C  , ,  �  #  �  �  W  �  W  #  �  #      C  , ,  �  �  �  5  W  5  W  �  �  �      C  , ,  �  �  �  �  W  �  W  �  �  �      C  , ,  �  [  �    W    W  [  �  [      C  , ,  �  �  �  m  W  m  W  �  �  �      C  , ,  �  +  �  �  W  �  W  +  �  +      C  , ,  �  �  �  =  W  =  W  �  �  �      C  , ,  �  �  �  �  W  �  W  �  �  �      C  , ,  �  c  �     W     W  c  �  c      C  , ,  �   �  �  !u  W  !u  W   �  �   �      C  , ,  �  "3  �  "�  W  "�  W  "3  �  "3      C  , ,  �  #�  �  $E  W  $E  W  #�  �  #�      C  , ,  �  %  �  %�  W  %�  W  %  �  %      C  , ,  �  &k  �  '  W  '  W  &k  �  &k      C  , ,  E  �  E  5  �  5  �  �  E  �      C  , ,  E  �  E  �  �  �  �  �  E  �      C  , ,  E  [  E    �    �  [  E  [      C  , ,  E  �  E  m  �  m  �  �  E  �      C  , ,  E  +  E  �  �  �  �  +  E  +      C  , ,  E  �  E  =  �  =  �  �  E  �      C  , ,  E  �  E  �  �  �  �  �  E  �      C  , ,  E  c  E     �     �  c  E  c      C  , ,  E   �  E  !u  �  !u  �   �  E   �      C  , ,  E  "3  E  "�  �  "�  �  "3  E  "3      C  , ,  �   s  �    �    �   s  �   s      C  , ,  �  �  �  �  �  �  �  �  �  �      C  , ,  �  C  �  �  �  �  �  C  �  C      C  , ,  �  �  �  U  �  U  �  �  �  �      C  , ,  �    �  �  �  �  �    �        C  , ,  �  {  �  %  �  %  �  {  �  {      C  , ,  �  �  �  	�  �  	�  �  �  �  �      C  , ,  �  
K  �  
�  �  
�  �  
K  �  
K      B  , ,   A  O3   A  O�   �  O�   �  O3   A  O3      B  , ,  �  O3  �  O�  S  O�  S  O3  �  O3      B  , ,    O3    O�  �  O�  �  O3    O3      B  , ,  �  O3  �  O�  �  O�  �  O3  �  O3      B  , ,  E  O3  E  O�  �  O�  �  O3  E  O3      B  , ,  �  O3  �  O�  W  O�  W  O3  �  O3      B  , ,  r  O3  r  O�    O�    O3  r  O3      B  , ,  �  O3  �  O�  �  O�  �  O3  �  O3      B  , ,  B  O3  B  O�  �  O�  �  O3  B  O3      B  , ,   A  v�   A  w=   �  w=   �  v�   A  v�      B  , ,  �  v�  �  w=  S  w=  S  v�  �  v�      B  , ,    v�    w=  �  w=  �  v�    v�      B  , ,  �  v�  �  w=  �  w=  �  v�  �  v�      B  , ,  E  v�  E  w=  �  w=  �  v�  E  v�      B  , ,  �  v�  �  w=  W  w=  W  v�  �  v�      B  , ,  r  v�  r  w=    w=    v�  r  v�      B  , ,  �  v�  �  w=  �  w=  �  v�  �  v�      B  , ,  B  v�  B  w=  �  w=  �  v�  B  v�      B  , ,  �  �C  �  ��  �  ��  �  �C  �  �C      B  , ,  E  �C  E  ��  �  ��  �  �C  E  �C      B  , ,  �  �C  �  ��  W  ��  W  �C  �  �C      B  , ,  r  �C  r  ��    ��    �C  r  �C      B  , ,  �  �C  �  ��  �  ��  �  �C  �  �C      B  , ,  B  �C  B  ��  �  ��  �  �C  B  �C      B  , ,  E  �K  E  ��  �  ��  �  �K  E  �K      B  , ,  E  ��  E  �]  �  �]  �  ��  E  ��      B  , ,  E  �  E  ��  �  ��  �  �  E  �      B  , ,  E  ��  E  �-  �  �-  �  ��  E  ��      B  , ,  E  ��  E  ��  �  ��  �  ��  E  ��      B  , ,  E  �S  E  ��  �  ��  �  �S  E  �S      B  , ,  E  ��  E  �e  �  �e  �  ��  E  ��      B  , ,  E  �#  E  ��  �  ��  �  �#  E  �#      B  , ,  E  ��  E  �U  �  �U  �  ��  E  ��      B  , ,  �  ��  �  �U  W  �U  W  ��  �  ��      B  , ,  �  �  �  ��  W  ��  W  �  �  �      B  , ,  �  �{  �  �%  W  �%  W  �{  �  �{      B  , ,  �  ��  �  ��  W  ��  W  ��  �  ��      B  , ,  �  �K  �  ��  W  ��  W  �K  �  �K      B  , ,  �  ��  �  �]  W  �]  W  ��  �  ��      B  , ,  �  �  �  ��  W  ��  W  �  �  �      B  , ,  �  ��  �  �-  W  �-  W  ��  �  ��      B  , ,  �  ��  �  ��  W  ��  W  ��  �  ��      B  , ,  �  �S  �  ��  W  ��  W  �S  �  �S      B  , ,  �  ��  �  �e  W  �e  W  ��  �  ��      B  , ,  �  �#  �  ��  W  ��  W  �#  �  �#      B  , ,  E  �  E  ��  �  ��  �  �  E  �      B  , ,  r  ��  r  �U    �U    ��  r  ��      B  , ,  r  �  r  ��    ��    �  r  �      B  , ,  r  �{  r  �%    �%    �{  r  �{      B  , ,  r  ��  r  ��    ��    ��  r  ��      B  , ,  r  �K  r  ��    ��    �K  r  �K      B  , ,  r  ��  r  �]    �]    ��  r  ��      B  , ,  r  �  r  ��    ��    �  r  �      B  , ,  r  ��  r  �-    �-    ��  r  ��      B  , ,  r  ��  r  ��    ��    ��  r  ��      B  , ,  r  �S  r  ��    ��    �S  r  �S      B  , ,  r  ��  r  �e    �e    ��  r  ��      B  , ,  r  �#  r  ��    ��    �#  r  �#      B  , ,  E  �{  E  �%  �  �%  �  �{  E  �{      B  , ,  �  ��  �  �U  �  �U  �  ��  �  ��      B  , ,  �  �  �  ��  �  ��  �  �  �  �      B  , ,  �  �{  �  �%  �  �%  �  �{  �  �{      B  , ,  �  ��  �  ��  �  ��  �  ��  �  ��      B  , ,  �  �K  �  ��  �  ��  �  �K  �  �K      B  , ,  �  ��  �  �]  �  �]  �  ��  �  ��      B  , ,  �  �  �  ��  �  ��  �  �  �  �      B  , ,  �  ��  �  �-  �  �-  �  ��  �  ��      B  , ,  �  ��  �  ��  �  ��  �  ��  �  ��      B  , ,  �  �S  �  ��  �  ��  �  �S  �  �S      B  , ,  �  ��  �  �e  �  �e  �  ��  �  ��      B  , ,  �  �#  �  ��  �  ��  �  �#  �  �#      B  , ,  E  ��  E  ��  �  ��  �  ��  E  ��      B  , ,  B  ��  B  �U  �  �U  �  ��  B  ��      B  , ,  B  �  B  ��  �  ��  �  �  B  �      B  , ,  B  �{  B  �%  �  �%  �  �{  B  �{      B  , ,  B  ��  B  ��  �  ��  �  ��  B  ��      B  , ,  B  �K  B  ��  �  ��  �  �K  B  �K      B  , ,  B  ��  B  �]  �  �]  �  ��  B  ��      B  , ,  B  �  B  ��  �  ��  �  �  B  �      B  , ,  B  ��  B  �-  �  �-  �  ��  B  ��      B  , ,  B  ��  B  ��  �  ��  �  ��  B  ��      B  , ,  B  �S  B  ��  �  ��  �  �S  B  �S      B  , ,  B  ��  B  �e  �  �e  �  ��  B  ��      B  , ,  B  �#  B  ��  �  ��  �  �#  B  �#      B  , ,  �  �S  �  ��  �  ��  �  �S  �  �S      B  , ,  �  ��  �  �e  �  �e  �  ��  �  ��      B  , ,  �  �#  �  ��  �  ��  �  �#  �  �#      B  , ,  �  ��  �  �U  �  �U  �  ��  �  ��      B  , ,  �  �  �  ��  �  ��  �  �  �  �      B  , ,  G  �X  G  �  �  �  �  �X  G  �X      B  , ,  �  �X  �  �  Y  �  Y  �X  �  �X      B  , ,    �X    �  �  �  �  �X    �X      B  , ,    �X    �  )  �  )  �X    �X      B  , ,  �  �{  �  �%  �  �%  �  �{  �  �{      B  , ,  �  ��  �  ��  �  ��  �  ��  �  ��      B  , ,  �  �K  �  ��  �  ��  �  �K  �  �K      B  , ,  �  ��  �  �]  �  �]  �  ��  �  ��      B  , ,  �  �  �  ��  �  ��  �  �  �  �      B  , ,  �  ��  �  �-  �  �-  �  ��  �  ��      B  , ,  �  ��  �  ��  �  ��  �  ��  �  ��      B  , ,  �  �k  �  �  �  �  �  �k  �  �k      B  , ,  �  ��  �  �}  �  �}  �  ��  �  ��      B  , ,  �  �;  �  ��  �  ��  �  �;  �  �;      B  , ,  �  ��  �  �M  �  �M  �  ��  �  ��      B  , ,  �  w�  �  x�  �  x�  �  w�  �  w�      B  , ,  �  �  �  ��  �  ��  �  �  �  �      B  , ,  �  �s  �  �  �  �  �  �s  �  �s      B  , ,  �  z�  �  {u  �  {u  �  z�  �  z�      B  , ,  �  ��  �  ��  �  ��  �  ��  �  ��      B  , ,  �    �  �  �  �  �    �        B  , ,  �  |3  �  |�  �  |�  �  |3  �  |3      B  , ,  �  yc  �  z  �  z  �  yc  �  yc      B  , ,  �  }�  �  ~E  �  ~E  �  }�  �  }�      B  , ,  �  ��  �  �}  W  �}  W  ��  �  ��      B  , ,  �  �;  �  ��  W  ��  W  �;  �  �;      B  , ,  �  ��  �  �M  W  �M  W  ��  �  ��      B  , ,  �  �  �  ��  W  ��  W  �  �  �      B  , ,  �  �s  �  �  W  �  W  �s  �  �s      B  , ,  �  ��  �  ��  W  ��  W  ��  �  ��      B  , ,  E  yc  E  z  �  z  �  yc  E  yc      B  , ,  E  z�  E  {u  �  {u  �  z�  E  z�      B  , ,  E  |3  E  |�  �  |�  �  |3  E  |3      B  , ,  E  }�  E  ~E  �  ~E  �  }�  E  }�      B  , ,  E    E  �  �  �  �    E        B  , ,  E  �k  E  �  �  �  �  �k  E  �k      B  , ,  �  w�  �  x�  �  x�  �  w�  �  w�      B  , ,  �  yc  �  z  �  z  �  yc  �  yc      B  , ,  �  z�  �  {u  �  {u  �  z�  �  z�      B  , ,  �  |3  �  |�  �  |�  �  |3  �  |3      B  , ,  �  }�  �  ~E  �  ~E  �  }�  �  }�      B  , ,  �    �  �  �  �  �    �        B  , ,  �  �k  �  �  �  �  �  �k  �  �k      B  , ,  �  ��  �  �}  �  �}  �  ��  �  ��      B  , ,  �  �;  �  ��  �  ��  �  �;  �  �;      B  , ,  �  ��  �  �M  �  �M  �  ��  �  ��      B  , ,  �  �  �  ��  �  ��  �  �  �  �      B  , ,  �  �s  �  �  �  �  �  �s  �  �s      B  , ,  �  ��  �  ��  �  ��  �  ��  �  ��      B  , ,  E  ��  E  �}  �  �}  �  ��  E  ��      B  , ,  E  �;  E  ��  �  ��  �  �;  E  �;      B  , ,  E  ��  E  �M  �  �M  �  ��  E  ��      B  , ,  E  �  E  ��  �  ��  �  �  E  �      B  , ,  E  �s  E  �  �  �  �  �s  E  �s      B  , ,  E  ��  E  ��  �  ��  �  ��  E  ��      B  , ,  E  w�  E  x�  �  x�  �  w�  E  w�      B  , ,  �  w�  �  x�  W  x�  W  w�  �  w�      B  , ,  �  yc  �  z  W  z  W  yc  �  yc      B  , ,  �  z�  �  {u  W  {u  W  z�  �  z�      B  , ,  �  |3  �  |�  W  |�  W  |3  �  |3      B  , ,  �  }�  �  ~E  W  ~E  W  }�  �  }�      B  , ,  r  w�  r  x�    x�    w�  r  w�      B  , ,  r  yc  r  z    z    yc  r  yc      B  , ,  B  w�  B  x�  �  x�  �  w�  B  w�      B  , ,  B  yc  B  z  �  z  �  yc  B  yc      B  , ,  B  z�  B  {u  �  {u  �  z�  B  z�      B  , ,  B  |3  B  |�  �  |�  �  |3  B  |3      B  , ,  B  }�  B  ~E  �  ~E  �  }�  B  }�      B  , ,  B    B  �  �  �  �    B        B  , ,  B  �k  B  �  �  �  �  �k  B  �k      B  , ,  B  ��  B  �}  �  �}  �  ��  B  ��      B  , ,  B  �;  B  ��  �  ��  �  �;  B  �;      B  , ,  B  ��  B  �M  �  �M  �  ��  B  ��      B  , ,  B  �  B  ��  �  ��  �  �  B  �      B  , ,  B  �s  B  �  �  �  �  �s  B  �s      B  , ,  B  ��  B  ��  �  ��  �  ��  B  ��      B  , ,  r  z�  r  {u    {u    z�  r  z�      B  , ,  r  |3  r  |�    |�    |3  r  |3      B  , ,  r  }�  r  ~E    ~E    }�  r  }�      B  , ,  r    r  �    �      r        B  , ,  r  �k  r  �    �    �k  r  �k      B  , ,  r  ��  r  �}    �}    ��  r  ��      B  , ,  r  �;  r  ��    ��    �;  r  �;      B  , ,  r  ��  r  �M    �M    ��  r  ��      B  , ,  r  �  r  ��    ��    �  r  �      B  , ,  r  �s  r  �    �    �s  r  �s      B  , ,  r  ��  r  ��    ��    ��  r  ��      B  , ,  �    �  �  W  �  W    �        B  , ,  �  �k  �  �  W  �  W  �k  �  �k      B  , ,   A     A  �   �  �   �     A        B  , ,   A  �k   A  �   �  �   �  �k   A  �k      B  , ,   A  ��   A  �}   �  �}   �  ��   A  ��      B  , ,   A  �;   A  ��   �  ��   �  �;   A  �;      B  , ,   A  ��   A  �M   �  �M   �  ��   A  ��      B  , ,   A  �   A  ��   �  ��   �  �   A  �      B  , ,   A  �s   A  �   �  �   �  �s   A  �s      B  , ,   A  ��   A  ��   �  ��   �  ��   A  ��      B  , ,   A  �C   A  ��   �  ��   �  �C   A  �C      B  , ,   A  ��   A  �U   �  �U   �  ��   A  ��      B  , ,   A  �   A  ��   �  ��   �  �   A  �      B  , ,   A  �{   A  �%   �  �%   �  �{   A  �{      B  , ,   A  ��   A  ��   �  ��   �  ��   A  ��      B  , ,   A  �K   A  ��   �  ��   �  �K   A  �K      B  , ,   A  ��   A  �]   �  �]   �  ��   A  ��      B  , ,   A  �   A  ��   �  ��   �  �   A  �      B  , ,   A  ��   A  �-   �  �-   �  ��   A  ��      B  , ,   A  ��   A  ��   �  ��   �  ��   A  ��      B  , ,   A  �S   A  ��   �  ��   �  �S   A  �S      B  , ,   A  ��   A  �e   �  �e   �  ��   A  ��      B  , ,   A  �#   A  ��   �  ��   �  �#   A  �#      B  , ,   A  w�   A  x�   �  x�   �  w�   A  w�      B  , ,  �  w�  �  x�  S  x�  S  w�  �  w�      B  , ,  �  yc  �  z  S  z  S  yc  �  yc      B  , ,  �  z�  �  {u  S  {u  S  z�  �  z�      B  , ,  �  |3  �  |�  S  |�  S  |3  �  |3      B  , ,  �  }�  �  ~E  S  ~E  S  }�  �  }�      B  , ,  �    �  �  S  �  S    �        B  , ,  �  �k  �  �  S  �  S  �k  �  �k      B  , ,  �  ��  �  �}  S  �}  S  ��  �  ��      B  , ,  �  �;  �  ��  S  ��  S  �;  �  �;      B  , ,  �  ��  �  �M  S  �M  S  ��  �  ��      B  , ,  �  �  �  ��  S  ��  S  �  �  �      B  , ,  �  �s  �  �  S  �  S  �s  �  �s      B  , ,  �  ��  �  ��  S  ��  S  ��  �  ��      B  , ,  �  �C  �  ��  S  ��  S  �C  �  �C      B  , ,  �  ��  �  �U  S  �U  S  ��  �  ��      B  , ,  �  �  �  ��  S  ��  S  �  �  �      B  , ,  �  �{  �  �%  S  �%  S  �{  �  �{      B  , ,  �  ��  �  ��  S  ��  S  ��  �  ��      B  , ,  �  �K  �  ��  S  ��  S  �K  �  �K      B  , ,  �  ��  �  �]  S  �]  S  ��  �  ��      B  , ,  �  �  �  ��  S  ��  S  �  �  �      B  , ,  �  ��  �  �-  S  �-  S  ��  �  ��      B  , ,  �  ��  �  ��  S  ��  S  ��  �  ��      B  , ,  �  �S  �  ��  S  ��  S  �S  �  �S      B  , ,  �  ��  �  �e  S  �e  S  ��  �  ��      B  , ,  �  �#  �  ��  S  ��  S  �#  �  �#      B  , ,   A  yc   A  z   �  z   �  yc   A  yc      B  , ,    w�    x�  �  x�  �  w�    w�      B  , ,    yc    z  �  z  �  yc    yc      B  , ,    z�    {u  �  {u  �  z�    z�      B  , ,    |3    |�  �  |�  �  |3    |3      B  , ,    }�    ~E  �  ~E  �  }�    }�      B  , ,        �  �  �  �            B  , ,    �k    �  �  �  �  �k    �k      B  , ,    ��    �}  �  �}  �  ��    ��      B  , ,    �;    ��  �  ��  �  �;    �;      B  , ,    ��    �M  �  �M  �  ��    ��      B  , ,    �    ��  �  ��  �  �    �      B  , ,    �s    �  �  �  �  �s    �s      B  , ,    ��    ��  �  ��  �  ��    ��      B  , ,    �C    ��  �  ��  �  �C    �C      B  , ,    ��    �U  �  �U  �  ��    ��      B  , ,    �    ��  �  ��  �  �    �      B  , ,    �{    �%  �  �%  �  �{    �{      B  , ,    ��    ��  �  ��  �  ��    ��      B  , ,    �K    ��  �  ��  �  �K    �K      B  , ,    ��    �]  �  �]  �  ��    ��      B  , ,    �    ��  �  ��  �  �    �      B  , ,    ��    �-  �  �-  �  ��    ��      B  , ,    ��    ��  �  ��  �  ��    ��      B  , ,    �S    ��  �  ��  �  �S    �S      B  , ,    ��    �e  �  �e  �  ��    ��      B  , ,    �#    ��  �  ��  �  �#    �#      B  , ,   A  z�   A  {u   �  {u   �  z�   A  z�      B  , ,   A  |3   A  |�   �  |�   �  |3   A  |3      B  , ,   A  }�   A  ~E   �  ~E   �  }�   A  }�      B  , ,  o  �X  o  �    �    �X  o  �X      B  , ,  �  �X  �  �  �  �  �  �X  �  �X      B  , ,  ?  �X  ?  �  �  �  �  �X  ?  �X      B  , ,  �  �X  �  �  	Q  �  	Q  �X  �  �X      B  , ,  
  �X  
  �  
�  �  
�  �X  
  �X      B  , ,  w  �X  w  �  !  �  !  �X  w  �X      B  , ,  �  �X  �  �  �  �  �  �X  �  �X      B  , ,  �  W�  �  XM  S  XM  S  W�  �  W�      B  , ,  �  Y  �  Y�  S  Y�  S  Y  �  Y      B  , ,   A  R   A  R�   �  R�   �  R   A  R      B  , ,    P�    QE  �  QE  �  P�    P�      B  , ,    R    R�  �  R�  �  R    R      B  , ,    Sk    T  �  T  �  Sk    Sk      B  , ,    T�    U}  �  U}  �  T�    T�      B  , ,    V;    V�  �  V�  �  V;    V;      B  , ,    W�    XM  �  XM  �  W�    W�      B  , ,   A  T�   A  U}   �  U}   �  T�   A  T�      B  , ,    Y    Y�  �  Y�  �  Y    Y      B  , ,    Zs    [  �  [  �  Zs    Zs      B  , ,    [�    \�  �  \�  �  [�    [�      B  , ,    ]C    ]�  �  ]�  �  ]C    ]C      B  , ,    ^�    _U  �  _U  �  ^�    ^�      B  , ,    `    `�  �  `�  �  `    `      B  , ,    a{    b%  �  b%  �  a{    a{      B  , ,    b�    c�  �  c�  �  b�    b�      B  , ,    dK    d�  �  d�  �  dK    dK      B  , ,    e�    f]  �  f]  �  e�    e�      B  , ,    g    g�  �  g�  �  g    g      B  , ,    h�    i-  �  i-  �  h�    h�      B  , ,    i�    j�  �  j�  �  i�    i�      B  , ,    kS    k�  �  k�  �  kS    kS      B  , ,    l�    me  �  me  �  l�    l�      B  , ,   A  Y   A  Y�   �  Y�   �  Y   A  Y      B  , ,    n#    n�  �  n�  �  n#    n#      B  , ,    o�    p5  �  p5  �  o�    o�      B  , ,    p�    q�  �  q�  �  p�    p�      B  , ,    r[    s  �  s  �  r[    r[      B  , ,    s�    tm  �  tm  �  s�    s�      B  , ,    u+    u�  �  u�  �  u+    u+      B  , ,  �  Zs  �  [  S  [  S  Zs  �  Zs      B  , ,  �  [�  �  \�  S  \�  S  [�  �  [�      B  , ,  �  ]C  �  ]�  S  ]�  S  ]C  �  ]C      B  , ,  �  ^�  �  _U  S  _U  S  ^�  �  ^�      B  , ,  �  `  �  `�  S  `�  S  `  �  `      B  , ,  �  a{  �  b%  S  b%  S  a{  �  a{      B  , ,   A  V;   A  V�   �  V�   �  V;   A  V;      B  , ,  �  b�  �  c�  S  c�  S  b�  �  b�      B  , ,  �  dK  �  d�  S  d�  S  dK  �  dK      B  , ,  �  e�  �  f]  S  f]  S  e�  �  e�      B  , ,  �  g  �  g�  S  g�  S  g  �  g      B  , ,  �  h�  �  i-  S  i-  S  h�  �  h�      B  , ,  �  i�  �  j�  S  j�  S  i�  �  i�      B  , ,  �  kS  �  k�  S  k�  S  kS  �  kS      B  , ,  �  l�  �  me  S  me  S  l�  �  l�      B  , ,  �  n#  �  n�  S  n�  S  n#  �  n#      B  , ,  �  o�  �  p5  S  p5  S  o�  �  o�      B  , ,  �  p�  �  q�  S  q�  S  p�  �  p�      B  , ,  �  r[  �  s  S  s  S  r[  �  r[      B  , ,  �  s�  �  tm  S  tm  S  s�  �  s�      B  , ,  �  u+  �  u�  S  u�  S  u+  �  u+      B  , ,   A  Zs   A  [   �  [   �  Zs   A  Zs      B  , ,   A  g   A  g�   �  g�   �  g   A  g      B  , ,   A  h�   A  i-   �  i-   �  h�   A  h�      B  , ,   A  i�   A  j�   �  j�   �  i�   A  i�      B  , ,   A  kS   A  k�   �  k�   �  kS   A  kS      B  , ,   A  l�   A  me   �  me   �  l�   A  l�      B  , ,   A  n#   A  n�   �  n�   �  n#   A  n#      B  , ,   A  o�   A  p5   �  p5   �  o�   A  o�      B  , ,   A  Sk   A  T   �  T   �  Sk   A  Sk      B  , ,   A  p�   A  q�   �  q�   �  p�   A  p�      B  , ,   A  r[   A  s   �  s   �  r[   A  r[      B  , ,   A  s�   A  tm   �  tm   �  s�   A  s�      B  , ,   A  u+   A  u�   �  u�   �  u+   A  u+      B  , ,   A  [�   A  \�   �  \�   �  [�   A  [�      B  , ,   A  ]C   A  ]�   �  ]�   �  ]C   A  ]C      B  , ,   A  ^�   A  _U   �  _U   �  ^�   A  ^�      B  , ,   A  `   A  `�   �  `�   �  `   A  `      B  , ,   A  a{   A  b%   �  b%   �  a{   A  a{      B  , ,   A  b�   A  c�   �  c�   �  b�   A  b�      B  , ,   A  dK   A  d�   �  d�   �  dK   A  dK      B  , ,   A  e�   A  f]   �  f]   �  e�   A  e�      B  , ,   A  P�   A  QE   �  QE   �  P�   A  P�      B  , ,  �  P�  �  QE  S  QE  S  P�  �  P�      B  , ,  �  R  �  R�  S  R�  S  R  �  R      B  , ,  �  Sk  �  T  S  T  S  Sk  �  Sk      B  , ,   A  W�   A  XM   �  XM   �  W�   A  W�      B  , ,  �  T�  �  U}  S  U}  S  T�  �  T�      B  , ,  �  V;  �  V�  S  V�  S  V;  �  V;      B  , ,  r  b�  r  c�    c�    b�  r  b�      B  , ,  �  b�  �  c�  �  c�  �  b�  �  b�      B  , ,  �  b�  �  c�  W  c�  W  b�  �  b�      B  , ,  E  b�  E  c�  �  c�  �  b�  E  b�      B  , ,  B  b�  B  c�  �  c�  �  b�  B  b�      B  , ,  �  b�  �  c�  �  c�  �  b�  �  b�      B  , ,  r  kS  r  k�    k�    kS  r  kS      B  , ,  r  l�  r  me    me    l�  r  l�      B  , ,  r  n#  r  n�    n�    n#  r  n#      B  , ,  r  o�  r  p5    p5    o�  r  o�      B  , ,  r  p�  r  q�    q�    p�  r  p�      B  , ,  r  r[  r  s    s    r[  r  r[      B  , ,  r  s�  r  tm    tm    s�  r  s�      B  , ,  r  u+  r  u�    u�    u+  r  u+      B  , ,  r  dK  r  d�    d�    dK  r  dK      B  , ,  �  dK  �  d�  �  d�  �  dK  �  dK      B  , ,  �  e�  �  f]  �  f]  �  e�  �  e�      B  , ,  �  g  �  g�  �  g�  �  g  �  g      B  , ,  �  h�  �  i-  �  i-  �  h�  �  h�      B  , ,  �  i�  �  j�  �  j�  �  i�  �  i�      B  , ,  �  kS  �  k�  �  k�  �  kS  �  kS      B  , ,  �  l�  �  me  �  me  �  l�  �  l�      B  , ,  �  n#  �  n�  �  n�  �  n#  �  n#      B  , ,  �  o�  �  p5  �  p5  �  o�  �  o�      B  , ,  �  p�  �  q�  �  q�  �  p�  �  p�      B  , ,  �  r[  �  s  �  s  �  r[  �  r[      B  , ,  �  s�  �  tm  �  tm  �  s�  �  s�      B  , ,  �  u+  �  u�  �  u�  �  u+  �  u+      B  , ,  r  e�  r  f]    f]    e�  r  e�      B  , ,  �  dK  �  d�  W  d�  W  dK  �  dK      B  , ,  �  e�  �  f]  W  f]  W  e�  �  e�      B  , ,  �  g  �  g�  W  g�  W  g  �  g      B  , ,  �  h�  �  i-  W  i-  W  h�  �  h�      B  , ,  �  i�  �  j�  W  j�  W  i�  �  i�      B  , ,  �  kS  �  k�  W  k�  W  kS  �  kS      B  , ,  �  l�  �  me  W  me  W  l�  �  l�      B  , ,  �  n#  �  n�  W  n�  W  n#  �  n#      B  , ,  �  o�  �  p5  W  p5  W  o�  �  o�      B  , ,  �  p�  �  q�  W  q�  W  p�  �  p�      B  , ,  �  r[  �  s  W  s  W  r[  �  r[      B  , ,  �  s�  �  tm  W  tm  W  s�  �  s�      B  , ,  �  u+  �  u�  W  u�  W  u+  �  u+      B  , ,  r  g  r  g�    g�    g  r  g      B  , ,  E  dK  E  d�  �  d�  �  dK  E  dK      B  , ,  r  h�  r  i-    i-    h�  r  h�      B  , ,  B  dK  B  d�  �  d�  �  dK  B  dK      B  , ,  B  e�  B  f]  �  f]  �  e�  B  e�      B  , ,  B  g  B  g�  �  g�  �  g  B  g      B  , ,  B  h�  B  i-  �  i-  �  h�  B  h�      B  , ,  B  i�  B  j�  �  j�  �  i�  B  i�      B  , ,  B  kS  B  k�  �  k�  �  kS  B  kS      B  , ,  B  l�  B  me  �  me  �  l�  B  l�      B  , ,  B  n#  B  n�  �  n�  �  n#  B  n#      B  , ,  B  o�  B  p5  �  p5  �  o�  B  o�      B  , ,  B  p�  B  q�  �  q�  �  p�  B  p�      B  , ,  B  r[  B  s  �  s  �  r[  B  r[      B  , ,  B  s�  B  tm  �  tm  �  s�  B  s�      B  , ,  B  u+  B  u�  �  u�  �  u+  B  u+      B  , ,  E  e�  E  f]  �  f]  �  e�  E  e�      B  , ,  E  g  E  g�  �  g�  �  g  E  g      B  , ,  E  h�  E  i-  �  i-  �  h�  E  h�      B  , ,  E  i�  E  j�  �  j�  �  i�  E  i�      B  , ,  E  kS  E  k�  �  k�  �  kS  E  kS      B  , ,  E  l�  E  me  �  me  �  l�  E  l�      B  , ,  E  n#  E  n�  �  n�  �  n#  E  n#      B  , ,  E  o�  E  p5  �  p5  �  o�  E  o�      B  , ,  E  p�  E  q�  �  q�  �  p�  E  p�      B  , ,  E  r[  E  s  �  s  �  r[  E  r[      B  , ,  E  s�  E  tm  �  tm  �  s�  E  s�      B  , ,  E  u+  E  u�  �  u�  �  u+  E  u+      B  , ,  r  i�  r  j�    j�    i�  r  i�      B  , ,  �  kS  �  k�  �  k�  �  kS  �  kS      B  , ,  �  l�  �  me  �  me  �  l�  �  l�      B  , ,  �  n#  �  n�  �  n�  �  n#  �  n#      B  , ,  �  o�  �  p5  �  p5  �  o�  �  o�      B  , ,  �  p�  �  q�  �  q�  �  p�  �  p�      B  , ,  �  r[  �  s  �  s  �  r[  �  r[      B  , ,  �  s�  �  tm  �  tm  �  s�  �  s�      B  , ,  �  u+  �  u�  �  u�  �  u+  �  u+      B  , ,  �  dK  �  d�  �  d�  �  dK  �  dK      B  , ,  �  e�  �  f]  �  f]  �  e�  �  e�      B  , ,  �  g  �  g�  �  g�  �  g  �  g      B  , ,  �  h�  �  i-  �  i-  �  h�  �  h�      B  , ,  �  i�  �  j�  �  j�  �  i�  �  i�      B  , ,  �  R  �  R�  �  R�  �  R  �  R      B  , ,  �  Sk  �  T  �  T  �  Sk  �  Sk      B  , ,  �  T�  �  U}  �  U}  �  T�  �  T�      B  , ,  �  V;  �  V�  �  V�  �  V;  �  V;      B  , ,  �  W�  �  XM  �  XM  �  W�  �  W�      B  , ,  �  Y  �  Y�  �  Y�  �  Y  �  Y      B  , ,  �  Zs  �  [  �  [  �  Zs  �  Zs      B  , ,  �  [�  �  \�  �  \�  �  [�  �  [�      B  , ,  �  ]C  �  ]�  �  ]�  �  ]C  �  ]C      B  , ,  �  ^�  �  _U  �  _U  �  ^�  �  ^�      B  , ,  �  `  �  `�  �  `�  �  `  �  `      B  , ,  �  a{  �  b%  �  b%  �  a{  �  a{      B  , ,  �  P�  �  QE  �  QE  �  P�  �  P�      B  , ,  E  V;  E  V�  �  V�  �  V;  E  V;      B  , ,  E  W�  E  XM  �  XM  �  W�  E  W�      B  , ,  E  Y  E  Y�  �  Y�  �  Y  E  Y      B  , ,  E  Zs  E  [  �  [  �  Zs  E  Zs      B  , ,  E  [�  E  \�  �  \�  �  [�  E  [�      B  , ,  E  ]C  E  ]�  �  ]�  �  ]C  E  ]C      B  , ,  E  ^�  E  _U  �  _U  �  ^�  E  ^�      B  , ,  E  `  E  `�  �  `�  �  `  E  `      B  , ,  E  a{  E  b%  �  b%  �  a{  E  a{      B  , ,  �  T�  �  U}  �  U}  �  T�  �  T�      B  , ,  �  V;  �  V�  �  V�  �  V;  �  V;      B  , ,  B  P�  B  QE  �  QE  �  P�  B  P�      B  , ,  B  R  B  R�  �  R�  �  R  B  R      B  , ,  B  Sk  B  T  �  T  �  Sk  B  Sk      B  , ,  B  T�  B  U}  �  U}  �  T�  B  T�      B  , ,  B  V;  B  V�  �  V�  �  V;  B  V;      B  , ,  B  W�  B  XM  �  XM  �  W�  B  W�      B  , ,  B  Y  B  Y�  �  Y�  �  Y  B  Y      B  , ,  B  Zs  B  [  �  [  �  Zs  B  Zs      B  , ,  B  [�  B  \�  �  \�  �  [�  B  [�      B  , ,  B  ]C  B  ]�  �  ]�  �  ]C  B  ]C      B  , ,  B  ^�  B  _U  �  _U  �  ^�  B  ^�      B  , ,  B  `  B  `�  �  `�  �  `  B  `      B  , ,  B  a{  B  b%  �  b%  �  a{  B  a{      B  , ,  �  W�  �  XM  �  XM  �  W�  �  W�      B  , ,  �  Y  �  Y�  �  Y�  �  Y  �  Y      B  , ,  �  Zs  �  [  �  [  �  Zs  �  Zs      B  , ,  �  [�  �  \�  �  \�  �  [�  �  [�      B  , ,  �  ]C  �  ]�  �  ]�  �  ]C  �  ]C      B  , ,  �  ^�  �  _U  �  _U  �  ^�  �  ^�      B  , ,  �  `  �  `�  �  `�  �  `  �  `      B  , ,  �  a{  �  b%  �  b%  �  a{  �  a{      B  , ,  r  [�  r  \�    \�    [�  r  [�      B  , ,  r  ]C  r  ]�    ]�    ]C  r  ]C      B  , ,  r  ^�  r  _U    _U    ^�  r  ^�      B  , ,  r  `  r  `�    `�    `  r  `      B  , ,  r  a{  r  b%    b%    a{  r  a{      B  , ,  r  Sk  r  T    T    Sk  r  Sk      B  , ,  r  T�  r  U}    U}    T�  r  T�      B  , ,  r  V;  r  V�    V�    V;  r  V;      B  , ,  r  W�  r  XM    XM    W�  r  W�      B  , ,  r  Y  r  Y�    Y�    Y  r  Y      B  , ,  r  Zs  r  [    [    Zs  r  Zs      B  , ,  E  P�  E  QE  �  QE  �  P�  E  P�      B  , ,  �  P�  �  QE  W  QE  W  P�  �  P�      B  , ,  �  R  �  R�  W  R�  W  R  �  R      B  , ,  �  Sk  �  T  W  T  W  Sk  �  Sk      B  , ,  �  T�  �  U}  W  U}  W  T�  �  T�      B  , ,  �  V;  �  V�  W  V�  W  V;  �  V;      B  , ,  �  W�  �  XM  W  XM  W  W�  �  W�      B  , ,  �  Y  �  Y�  W  Y�  W  Y  �  Y      B  , ,  �  Zs  �  [  W  [  W  Zs  �  Zs      B  , ,  �  [�  �  \�  W  \�  W  [�  �  [�      B  , ,  �  ]C  �  ]�  W  ]�  W  ]C  �  ]C      B  , ,  �  ^�  �  _U  W  _U  W  ^�  �  ^�      B  , ,  �  `  �  `�  W  `�  W  `  �  `      B  , ,  �  a{  �  b%  W  b%  W  a{  �  a{      B  , ,  �  P�  �  QE  �  QE  �  P�  �  P�      B  , ,  �  R  �  R�  �  R�  �  R  �  R      B  , ,  �  Sk  �  T  �  T  �  Sk  �  Sk      B  , ,  E  R  E  R�  �  R�  �  R  E  R      B  , ,  E  Sk  E  T  �  T  �  Sk  E  Sk      B  , ,  E  T�  E  U}  �  U}  �  T�  E  T�      B  , ,  r  P�  r  QE    QE    P�  r  P�      B  , ,  r  R  r  R�    R�    R  r  R      B  , ,    '�    (}  �  (}  �  '�    '�      B  , ,  �  '�  �  (}  W  (}  W  '�  �  '�      B  , ,  �  '�  �  (}  S  (}  S  '�  �  '�      B  , ,  r  '�  r  (}    (}    '�  r  '�      B  , ,  �  '�  �  (}  �  (}  �  '�  �  '�      B  , ,  �  '�  �  (}  �  (}  �  '�  �  '�      B  , ,   A  '�   A  (}   �  (}   �  '�   A  '�      B  , ,  B  '�  B  (}  �  (}  �  '�  B  '�      B  , ,  E  '�  E  (}  �  (}  �  '�  E  '�      B  , ,  �  ;�  �  <-  W  <-  W  ;�  �  ;�      B  , ,  r  ;�  r  <-    <-    ;�  r  ;�      B  , ,  �  ;�  �  <-  �  <-  �  ;�  �  ;�      B  , ,  �  ;�  �  <-  �  <-  �  ;�  �  ;�      B  , ,  B  ;�  B  <-  �  <-  �  ;�  B  ;�      B  , ,  E  ;�  E  <-  �  <-  �  ;�  E  ;�      B  , ,  �  C�  �  D�  W  D�  W  C�  �  C�      B  , ,  �  E[  �  F  W  F  W  E[  �  E[      B  , ,  �  F�  �  Gm  W  Gm  W  F�  �  F�      B  , ,  �  H+  �  H�  W  H�  W  H+  �  H+      B  , ,  �  I�  �  J=  W  J=  W  I�  �  I�      B  , ,  �  J�  �  K�  W  K�  W  J�  �  J�      B  , ,  �  Lc  �  M  W  M  W  Lc  �  Lc      B  , ,  �  M�  �  Nu  W  Nu  W  M�  �  M�      B  , ,  �  <�  �  =�  W  =�  W  <�  �  <�      B  , ,  r  <�  r  =�    =�    <�  r  <�      B  , ,  r  >S  r  >�    >�    >S  r  >S      B  , ,  r  ?�  r  @e    @e    ?�  r  ?�      B  , ,  r  A#  r  A�    A�    A#  r  A#      B  , ,  r  B�  r  C5    C5    B�  r  B�      B  , ,  r  C�  r  D�    D�    C�  r  C�      B  , ,  r  E[  r  F    F    E[  r  E[      B  , ,  r  F�  r  Gm    Gm    F�  r  F�      B  , ,  r  H+  r  H�    H�    H+  r  H+      B  , ,  r  I�  r  J=    J=    I�  r  I�      B  , ,  r  J�  r  K�    K�    J�  r  J�      B  , ,  r  Lc  r  M    M    Lc  r  Lc      B  , ,  r  M�  r  Nu    Nu    M�  r  M�      B  , ,  �  >S  �  >�  W  >�  W  >S  �  >S      B  , ,  �  ?�  �  @e  W  @e  W  ?�  �  ?�      B  , ,  �  <�  �  =�  �  =�  �  <�  �  <�      B  , ,  �  >S  �  >�  �  >�  �  >S  �  >S      B  , ,  �  ?�  �  @e  �  @e  �  ?�  �  ?�      B  , ,  �  A#  �  A�  �  A�  �  A#  �  A#      B  , ,  �  B�  �  C5  �  C5  �  B�  �  B�      B  , ,  �  C�  �  D�  �  D�  �  C�  �  C�      B  , ,  �  E[  �  F  �  F  �  E[  �  E[      B  , ,  �  F�  �  Gm  �  Gm  �  F�  �  F�      B  , ,  �  H+  �  H�  �  H�  �  H+  �  H+      B  , ,  �  I�  �  J=  �  J=  �  I�  �  I�      B  , ,  �  J�  �  K�  �  K�  �  J�  �  J�      B  , ,  �  Lc  �  M  �  M  �  Lc  �  Lc      B  , ,  �  M�  �  Nu  �  Nu  �  M�  �  M�      B  , ,  �  A#  �  A�  W  A�  W  A#  �  A#      B  , ,  B  <�  B  =�  �  =�  �  <�  B  <�      B  , ,  B  >S  B  >�  �  >�  �  >S  B  >S      B  , ,  B  ?�  B  @e  �  @e  �  ?�  B  ?�      B  , ,  B  A#  B  A�  �  A�  �  A#  B  A#      B  , ,  B  B�  B  C5  �  C5  �  B�  B  B�      B  , ,  B  C�  B  D�  �  D�  �  C�  B  C�      B  , ,  B  E[  B  F  �  F  �  E[  B  E[      B  , ,  B  F�  B  Gm  �  Gm  �  F�  B  F�      B  , ,  B  H+  B  H�  �  H�  �  H+  B  H+      B  , ,  B  I�  B  J=  �  J=  �  I�  B  I�      B  , ,  B  J�  B  K�  �  K�  �  J�  B  J�      B  , ,  B  Lc  B  M  �  M  �  Lc  B  Lc      B  , ,  B  M�  B  Nu  �  Nu  �  M�  B  M�      B  , ,  �  B�  �  C5  W  C5  W  B�  �  B�      B  , ,  E  <�  E  =�  �  =�  �  <�  E  <�      B  , ,  E  >S  E  >�  �  >�  �  >S  E  >S      B  , ,  E  ?�  E  @e  �  @e  �  ?�  E  ?�      B  , ,  E  A#  E  A�  �  A�  �  A#  E  A#      B  , ,  E  B�  E  C5  �  C5  �  B�  E  B�      B  , ,  E  C�  E  D�  �  D�  �  C�  E  C�      B  , ,  E  E[  E  F  �  F  �  E[  E  E[      B  , ,  E  F�  E  Gm  �  Gm  �  F�  E  F�      B  , ,  E  H+  E  H�  �  H�  �  H+  E  H+      B  , ,  E  I�  E  J=  �  J=  �  I�  E  I�      B  , ,  E  J�  E  K�  �  K�  �  J�  E  J�      B  , ,  E  Lc  E  M  �  M  �  Lc  E  Lc      B  , ,  E  M�  E  Nu  �  Nu  �  M�  E  M�      B  , ,  �  A#  �  A�  �  A�  �  A#  �  A#      B  , ,  �  B�  �  C5  �  C5  �  B�  �  B�      B  , ,  �  C�  �  D�  �  D�  �  C�  �  C�      B  , ,  �  E[  �  F  �  F  �  E[  �  E[      B  , ,  �  F�  �  Gm  �  Gm  �  F�  �  F�      B  , ,  �  H+  �  H�  �  H�  �  H+  �  H+      B  , ,  �  I�  �  J=  �  J=  �  I�  �  I�      B  , ,  �  J�  �  K�  �  K�  �  J�  �  J�      B  , ,  �  Lc  �  M  �  M  �  Lc  �  Lc      B  , ,  �  M�  �  Nu  �  Nu  �  M�  �  M�      B  , ,  �  <�  �  =�  �  =�  �  <�  �  <�      B  , ,  �  >S  �  >�  �  >�  �  >S  �  >S      B  , ,  �  ?�  �  @e  �  @e  �  ?�  �  ?�      B  , ,  �  .�  �  /�  �  /�  �  .�  �  .�      B  , ,  �  0C  �  0�  �  0�  �  0C  �  0C      B  , ,  �  1�  �  2U  �  2U  �  1�  �  1�      B  , ,  �  3  �  3�  �  3�  �  3  �  3      B  , ,  �  4{  �  5%  �  5%  �  4{  �  4{      B  , ,  �  5�  �  6�  �  6�  �  5�  �  5�      B  , ,  �  7K  �  7�  �  7�  �  7K  �  7K      B  , ,  �  8�  �  9]  �  9]  �  8�  �  8�      B  , ,  �  :  �  :�  �  :�  �  :  �  :      B  , ,  �  );  �  )�  �  )�  �  );  �  );      B  , ,  �  *�  �  +M  �  +M  �  *�  �  *�      B  , ,  �  ,  �  ,�  �  ,�  �  ,  �  ,      B  , ,  �  -s  �  .  �  .  �  -s  �  -s      B  , ,  �  3  �  3�  W  3�  W  3  �  3      B  , ,  �  4{  �  5%  W  5%  W  4{  �  4{      B  , ,  �  );  �  )�  W  )�  W  );  �  );      B  , ,  �  *�  �  +M  W  +M  W  *�  �  *�      B  , ,  r  );  r  )�    )�    );  r  );      B  , ,  r  *�  r  +M    +M    *�  r  *�      B  , ,  r  ,  r  ,�    ,�    ,  r  ,      B  , ,  r  -s  r  .    .    -s  r  -s      B  , ,  �  .�  �  /�  W  /�  W  .�  �  .�      B  , ,  �  0C  �  0�  W  0�  W  0C  �  0C      B  , ,  B  );  B  )�  �  )�  �  );  B  );      B  , ,  B  *�  B  +M  �  +M  �  *�  B  *�      B  , ,  B  ,  B  ,�  �  ,�  �  ,  B  ,      B  , ,  B  -s  B  .  �  .  �  -s  B  -s      B  , ,  B  .�  B  /�  �  /�  �  .�  B  .�      B  , ,  B  0C  B  0�  �  0�  �  0C  B  0C      B  , ,  B  1�  B  2U  �  2U  �  1�  B  1�      B  , ,  B  3  B  3�  �  3�  �  3  B  3      B  , ,  B  4{  B  5%  �  5%  �  4{  B  4{      B  , ,  B  5�  B  6�  �  6�  �  5�  B  5�      B  , ,  B  7K  B  7�  �  7�  �  7K  B  7K      B  , ,  B  8�  B  9]  �  9]  �  8�  B  8�      B  , ,  B  :  B  :�  �  :�  �  :  B  :      B  , ,  r  .�  r  /�    /�    .�  r  .�      B  , ,  r  0C  r  0�    0�    0C  r  0C      B  , ,  �  ,  �  ,�  W  ,�  W  ,  �  ,      B  , ,  r  1�  r  2U    2U    1�  r  1�      B  , ,  r  3  r  3�    3�    3  r  3      B  , ,  r  4{  r  5%    5%    4{  r  4{      B  , ,  r  5�  r  6�    6�    5�  r  5�      B  , ,  r  7K  r  7�    7�    7K  r  7K      B  , ,  �  -s  �  .  W  .  W  -s  �  -s      B  , ,  �  );  �  )�  �  )�  �  );  �  );      B  , ,  �  *�  �  +M  �  +M  �  *�  �  *�      B  , ,  �  ,  �  ,�  �  ,�  �  ,  �  ,      B  , ,  �  -s  �  .  �  .  �  -s  �  -s      B  , ,  �  .�  �  /�  �  /�  �  .�  �  .�      B  , ,  �  1�  �  2U  W  2U  W  1�  �  1�      B  , ,  E  );  E  )�  �  )�  �  );  E  );      B  , ,  E  *�  E  +M  �  +M  �  *�  E  *�      B  , ,  E  ,  E  ,�  �  ,�  �  ,  E  ,      B  , ,  E  -s  E  .  �  .  �  -s  E  -s      B  , ,  E  .�  E  /�  �  /�  �  .�  E  .�      B  , ,  E  0C  E  0�  �  0�  �  0C  E  0C      B  , ,  E  1�  E  2U  �  2U  �  1�  E  1�      B  , ,  E  3  E  3�  �  3�  �  3  E  3      B  , ,  E  4{  E  5%  �  5%  �  4{  E  4{      B  , ,  E  5�  E  6�  �  6�  �  5�  E  5�      B  , ,  E  7K  E  7�  �  7�  �  7K  E  7K      B  , ,  E  8�  E  9]  �  9]  �  8�  E  8�      B  , ,  E  :  E  :�  �  :�  �  :  E  :      B  , ,  �  0C  �  0�  �  0�  �  0C  �  0C      B  , ,  �  1�  �  2U  �  2U  �  1�  �  1�      B  , ,  �  3  �  3�  �  3�  �  3  �  3      B  , ,  �  4{  �  5%  �  5%  �  4{  �  4{      B  , ,  �  5�  �  6�  �  6�  �  5�  �  5�      B  , ,  �  7K  �  7�  �  7�  �  7K  �  7K      B  , ,  �  8�  �  9]  �  9]  �  8�  �  8�      B  , ,  �  :  �  :�  �  :�  �  :  �  :      B  , ,  r  8�  r  9]    9]    8�  r  8�      B  , ,  r  :  r  :�    :�    :  r  :      B  , ,  �  5�  �  6�  W  6�  W  5�  �  5�      B  , ,  �  7K  �  7�  W  7�  W  7K  �  7K      B  , ,  �  8�  �  9]  W  9]  W  8�  �  8�      B  , ,  �  :  �  :�  W  :�  W  :  �  :      B  , ,   A  );   A  )�   �  )�   �  );   A  );      B  , ,   A  *�   A  +M   �  +M   �  *�   A  *�      B  , ,   A  ,   A  ,�   �  ,�   �  ,   A  ,      B  , ,   A  -s   A  .   �  .   �  -s   A  -s      B  , ,   A  .�   A  /�   �  /�   �  .�   A  .�      B  , ,   A  0C   A  0�   �  0�   �  0C   A  0C      B  , ,   A  1�   A  2U   �  2U   �  1�   A  1�      B  , ,   A  3   A  3�   �  3�   �  3   A  3      B  , ,   A  4{   A  5%   �  5%   �  4{   A  4{      B  , ,   A  5�   A  6�   �  6�   �  5�   A  5�      B  , ,   A  7K   A  7�   �  7�   �  7K   A  7K      B  , ,   A  8�   A  9]   �  9]   �  8�   A  8�      B  , ,   A  :   A  :�   �  :�   �  :   A  :      B  , ,   A  ;�   A  <-   �  <-   �  ;�   A  ;�      B  , ,   A  <�   A  =�   �  =�   �  <�   A  <�      B  , ,   A  >S   A  >�   �  >�   �  >S   A  >S      B  , ,   A  ?�   A  @e   �  @e   �  ?�   A  ?�      B  , ,   A  A#   A  A�   �  A�   �  A#   A  A#      B  , ,   A  B�   A  C5   �  C5   �  B�   A  B�      B  , ,   A  C�   A  D�   �  D�   �  C�   A  C�      B  , ,   A  E[   A  F   �  F   �  E[   A  E[      B  , ,   A  F�   A  Gm   �  Gm   �  F�   A  F�      B  , ,   A  H+   A  H�   �  H�   �  H+   A  H+      B  , ,  �  .�  �  /�  S  /�  S  .�  �  .�      B  , ,  �  0C  �  0�  S  0�  S  0C  �  0C      B  , ,  �  1�  �  2U  S  2U  S  1�  �  1�      B  , ,  �  3  �  3�  S  3�  S  3  �  3      B  , ,  �  4{  �  5%  S  5%  S  4{  �  4{      B  , ,  �  5�  �  6�  S  6�  S  5�  �  5�      B  , ,  �  7K  �  7�  S  7�  S  7K  �  7K      B  , ,  �  8�  �  9]  S  9]  S  8�  �  8�      B  , ,  �  :  �  :�  S  :�  S  :  �  :      B  , ,  �  ;�  �  <-  S  <-  S  ;�  �  ;�      B  , ,  �  <�  �  =�  S  =�  S  <�  �  <�      B  , ,  �  >S  �  >�  S  >�  S  >S  �  >S      B  , ,  �  ?�  �  @e  S  @e  S  ?�  �  ?�      B  , ,  �  A#  �  A�  S  A�  S  A#  �  A#      B  , ,  �  B�  �  C5  S  C5  S  B�  �  B�      B  , ,  �  C�  �  D�  S  D�  S  C�  �  C�      B  , ,  �  E[  �  F  S  F  S  E[  �  E[      B  , ,  �  F�  �  Gm  S  Gm  S  F�  �  F�      B  , ,  �  H+  �  H�  S  H�  S  H+  �  H+      B  , ,  �  I�  �  J=  S  J=  S  I�  �  I�      B  , ,  �  J�  �  K�  S  K�  S  J�  �  J�      B  , ,    0C    0�  �  0�  �  0C    0C      B  , ,    1�    2U  �  2U  �  1�    1�      B  , ,    3    3�  �  3�  �  3    3      B  , ,  �  Lc  �  M  S  M  S  Lc  �  Lc      B  , ,  �  M�  �  Nu  S  Nu  S  M�  �  M�      B  , ,   A  M�   A  Nu   �  Nu   �  M�   A  M�      B  , ,    4{    5%  �  5%  �  4{    4{      B  , ,    5�    6�  �  6�  �  5�    5�      B  , ,    7K    7�  �  7�  �  7K    7K      B  , ,    8�    9]  �  9]  �  8�    8�      B  , ,    :    :�  �  :�  �  :    :      B  , ,    ;�    <-  �  <-  �  ;�    ;�      B  , ,    <�    =�  �  =�  �  <�    <�      B  , ,    >S    >�  �  >�  �  >S    >S      B  , ,    ?�    @e  �  @e  �  ?�    ?�      B  , ,    A#    A�  �  A�  �  A#    A#      B  , ,    B�    C5  �  C5  �  B�    B�      B  , ,    C�    D�  �  D�  �  C�    C�      B  , ,    E[    F  �  F  �  E[    E[      B  , ,    F�    Gm  �  Gm  �  F�    F�      B  , ,    H+    H�  �  H�  �  H+    H+      B  , ,    I�    J=  �  J=  �  I�    I�      B  , ,    );    )�  �  )�  �  );    );      B  , ,    *�    +M  �  +M  �  *�    *�      B  , ,    ,    ,�  �  ,�  �  ,    ,      B  , ,    -s    .  �  .  �  -s    -s      B  , ,    J�    K�  �  K�  �  J�    J�      B  , ,    Lc    M  �  M  �  Lc    Lc      B  , ,    M�    Nu  �  Nu  �  M�    M�      B  , ,   A  Lc   A  M   �  M   �  Lc   A  Lc      B  , ,    .�    /�  �  /�  �  .�    .�      B  , ,  �  );  �  )�  S  )�  S  );  �  );      B  , ,  �  *�  �  +M  S  +M  S  *�  �  *�      B  , ,  �  ,  �  ,�  S  ,�  S  ,  �  ,      B  , ,  �  -s  �  .  S  .  S  -s  �  -s      B  , ,   A  I�   A  J=   �  J=   �  I�   A  I�      B  , ,   A  J�   A  K�   �  K�   �  J�   A  J�      B  , ,    "3    "�  �  "�  �  "3    "3      B  , ,    #�    $E  �  $E  �  #�    #�      B  , ,    %    %�  �  %�  �  %    %      B  , ,    &k    '  �  '  �  &k    &k      B  , ,        �  �  �  �            B  , ,    {    %  �  %  �  {    {      B  , ,    �    	�  �  	�  �  �    �      B  , ,    
K    
�  �  
�  �  
K    
K      B  , ,    �    ]  �  ]  �  �    �      B  , ,        �  �  �  �            B  , ,    �    -  �  -  �  �    �      B  , ,    �    �  �  �  �  �    �      B  , ,    S    �  �  �  �  S    S      B  , ,  �   s  �    S    S   s  �   s      B  , ,  �  �  �  �  S  �  S  �  �  �      B  , ,  �  C  �  �  S  �  S  C  �  C      B  , ,  �  �  �  U  S  U  S  �  �  �      B  , ,  �    �  �  S  �  S    �        B  , ,  �  {  �  %  S  %  S  {  �  {      B  , ,  �  �  �  	�  S  	�  S  �  �  �      B  , ,  �  
K  �  
�  S  
�  S  
K  �  
K      B  , ,  �  �  �  ]  S  ]  S  �  �  �      B  , ,   A   s   A     �     �   s   A   s      B  , ,   A  �   A  �   �  �   �  �   A  �      B  , ,   A  C   A  �   �  �   �  C   A  C      B  , ,   A  �   A  U   �  U   �  �   A  �      B  , ,  �    �  �  S  �  S    �        B  , ,  �  �  �  -  S  -  S  �  �  �      B  , ,  �  �  �  �  S  �  S  �  �  �      B  , ,  �  S  �  �  S  �  S  S  �  S      B  , ,  �  �  �  e  S  e  S  �  �  �      B  , ,  �  #  �  �  S  �  S  #  �  #      B  , ,  �  �  �  5  S  5  S  �  �  �      B  , ,  �  �  �  �  S  �  S  �  �  �      B  , ,  �  [  �    S    S  [  �  [      B  , ,  �  �  �  m  S  m  S  �  �  �      B  , ,  �  +  �  �  S  �  S  +  �  +      B  , ,  �  �  �  =  S  =  S  �  �  �      B  , ,  �  �  �  �  S  �  S  �  �  �      B  , ,  �  c  �     S     S  c  �  c      B  , ,  �   �  �  !u  S  !u  S   �  �   �      B  , ,  �  "3  �  "�  S  "�  S  "3  �  "3      B  , ,  �  #�  �  $E  S  $E  S  #�  �  #�      B  , ,  �  %  �  %�  S  %�  S  %  �  %      B  , ,  �  &k  �  '  S  '  S  &k  �  &k      B  , ,    �    e  �  e  �  �    �      B  , ,    #    �  �  �  �  #    #      B  , ,    �    5  �  5  �  �    �      B  , ,    �    �  �  �  �  �    �      B  , ,    [      �    �  [    [      B  , ,    �    m  �  m  �  �    �      B  , ,    +    �  �  �  �  +    +      B  , ,    �    =  �  =  �  �    �      B  , ,    �    �  �  �  �  �    �      B  , ,   A     A  �   �  �   �     A        B  , ,   A  {   A  %   �  %   �  {   A  {      B  , ,   A  �   A  	�   �  	�   �  �   A  �      B  , ,   A  
K   A  
�   �  
�   �  
K   A  
K      B  , ,   A  �   A  ]   �  ]   �  �   A  �      B  , ,   A     A  �   �  �   �     A        B  , ,   A  �   A  -   �  -   �  �   A  �      B  , ,   A  �   A  �   �  �   �  �   A  �      B  , ,   A  S   A  �   �  �   �  S   A  S      B  , ,   A  �   A  e   �  e   �  �   A  �      B  , ,   A  #   A  �   �  �   �  #   A  #      B  , ,   A  �   A  5   �  5   �  �   A  �      B  , ,   A  �   A  �   �  �   �  �   A  �      B  , ,   A  [   A     �     �  [   A  [      B  , ,   A  �   A  m   �  m   �  �   A  �      B  , ,   A  +   A  �   �  �   �  +   A  +      B  , ,   A  �   A  =   �  =   �  �   A  �      B  , ,   A  �   A  �   �  �   �  �   A  �      B  , ,   A  c   A      �      �  c   A  c      B  , ,   A   �   A  !u   �  !u   �   �   A   �      B  , ,   A  "3   A  "�   �  "�   �  "3   A  "3      B  , ,   A  #�   A  $E   �  $E   �  #�   A  #�      B  , ,   A  %   A  %�   �  %�   �  %   A  %      B  , ,   A  &k   A  '   �  '   �  &k   A  &k      B  , ,    c       �     �  c    c      B  , ,     �    !u  �  !u  �   �     �      B  , ,     s      �    �   s     s      B  , ,    �    �  �  �  �  �    �      B  , ,    C    �  �  �  �  C    C      B  , ,    �    U  �  U  �  �    �      B  , ,  �  #  �  �  �  �  �  #  �  #      B  , ,  r  #  r  �    �    #  r  #      B  , ,  B  #  B  �  �  �  �  #  B  #      B  , ,  �  #  �  �  �  �  �  #  �  #      B  , ,  E  #  E  �  �  �  �  #  E  #      B  , ,  �  #  �  �  W  �  W  #  �  #      B  , ,  r  �  r  m    m    �  r  �      B  , ,  �  &k  �  '  W  '  W  &k  �  &k      B  , ,  B  �  B  5  �  5  �  �  B  �      B  , ,  B  �  B  �  �  �  �  �  B  �      B  , ,  B  [  B    �    �  [  B  [      B  , ,  B  �  B  m  �  m  �  �  B  �      B  , ,  B  +  B  �  �  �  �  +  B  +      B  , ,  B  �  B  =  �  =  �  �  B  �      B  , ,  B  �  B  �  �  �  �  �  B  �      B  , ,  B  c  B     �     �  c  B  c      B  , ,  B   �  B  !u  �  !u  �   �  B   �      B  , ,  B  "3  B  "�  �  "�  �  "3  B  "3      B  , ,  B  #�  B  $E  �  $E  �  #�  B  #�      B  , ,  B  %  B  %�  �  %�  �  %  B  %      B  , ,  B  &k  B  '  �  '  �  &k  B  &k      B  , ,  r  +  r  �    �    +  r  +      B  , ,  r  �  r  =    =    �  r  �      B  , ,  r  �  r  �    �    �  r  �      B  , ,  r  c  r            c  r  c      B  , ,  r   �  r  !u    !u     �  r   �      B  , ,  r  "3  r  "�    "�    "3  r  "3      B  , ,  r  #�  r  $E    $E    #�  r  #�      B  , ,  r  %  r  %�    %�    %  r  %      B  , ,  r  �  r  5    5    �  r  �      B  , ,  �  �  �  5  �  5  �  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  �  [  �    �    �  [  �  [      B  , ,  �  �  �  m  �  m  �  �  �  �      B  , ,  �  +  �  �  �  �  �  +  �  +      B  , ,  r  �  r  �    �    �  r  �      B  , ,  E  �  E  5  �  5  �  �  E  �      B  , ,  E  �  E  �  �  �  �  �  E  �      B  , ,  E  [  E    �    �  [  E  [      B  , ,  E  �  E  m  �  m  �  �  E  �      B  , ,  E  +  E  �  �  �  �  +  E  +      B  , ,  E  �  E  =  �  =  �  �  E  �      B  , ,  E  �  E  �  �  �  �  �  E  �      B  , ,  E  c  E     �     �  c  E  c      B  , ,  E   �  E  !u  �  !u  �   �  E   �      B  , ,  E  "3  E  "�  �  "�  �  "3  E  "3      B  , ,  E  #�  E  $E  �  $E  �  #�  E  #�      B  , ,  E  %  E  %�  �  %�  �  %  E  %      B  , ,  E  &k  E  '  �  '  �  &k  E  &k      B  , ,  �  �  �  =  �  =  �  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  �  c  �     �     �  c  �  c      B  , ,  �   �  �  !u  �  !u  �   �  �   �      B  , ,  �  "3  �  "�  �  "�  �  "3  �  "3      B  , ,  �  #�  �  $E  �  $E  �  #�  �  #�      B  , ,  �  %  �  %�  �  %�  �  %  �  %      B  , ,  �  &k  �  '  �  '  �  &k  �  &k      B  , ,  r  &k  r  '    '    &k  r  &k      B  , ,  r  [  r          [  r  [      B  , ,  �  �  �  5  W  5  W  �  �  �      B  , ,  �  �  �  �  W  �  W  �  �  �      B  , ,  �  [  �    W    W  [  �  [      B  , ,  �  �  �  m  W  m  W  �  �  �      B  , ,  �  +  �  �  W  �  W  +  �  +      B  , ,  �  �  �  =  W  =  W  �  �  �      B  , ,  �  �  �  �  W  �  W  �  �  �      B  , ,  �  c  �     W     W  c  �  c      B  , ,  �   �  �  !u  W  !u  W   �  �   �      B  , ,  �  "3  �  "�  W  "�  W  "3  �  "3      B  , ,  �  #�  �  $E  W  $E  W  #�  �  #�      B  , ,  �  %  �  %�  W  %�  W  %  �  %      B  , ,  �  +  �  �  �  �  �  +  �  +      B  , ,  �  �  �  =  �  =  �  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  �  c  �     �     �  c  �  c      B  , ,  �   �  �  !u  �  !u  �   �  �   �      B  , ,  �  "3  �  "�  �  "�  �  "3  �  "3      B  , ,  �  #�  �  $E  �  $E  �  #�  �  #�      B  , ,  �  %  �  %�  �  %�  �  %  �  %      B  , ,  �  &k  �  '  �  '  �  &k  �  &k      B  , ,  �  �  �  5  �  5  �  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  �  [  �    �    �  [  �  [      B  , ,  �  �  �  m  �  m  �  �  �  �      B  , ,  �  
K  �  
�  �  
�  �  
K  �  
K      B  , ,  �  �  �  -  �  -  �  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  �  S  �  �  �  �  �  S  �  S      B  , ,  �  �  �  e  �  e  �  �  �  �      B  , ,  �  �  �  ]  �  ]  �  �  �  �      B  , ,  �    �  �  �  �  �    �        B  , ,  �   s  �    �    �   s  �   s      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  �  C  �  �  �  �  �  C  �  C      B  , ,  �  �  �  U  �  U  �  �  �  �      B  , ,  �    �  �  �  �  �    �        B  , ,  �  {  �  %  �  %  �  {  �  {      B  , ,  �  �  �  	�  �  	�  �  �  �  �      B  , ,  �  {  �  %  �  %  �  {  �  {      B  , ,  �  �  �  	�  �  	�  �  �  �  �      B  , ,  �  
K  �  
�  �  
�  �  
K  �  
K      B  , ,  �  �  �  ]  �  ]  �  �  �  �      B  , ,  �    �  �  �  �  �    �        B  , ,  �  �  �  -  �  -  �  �  �  �      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  �  S  �  �  �  �  �  S  �  S      B  , ,  �  �  �  e  �  e  �  �  �  �      B  , ,  E  �  E  	�  �  	�  �  �  E  �      B  , ,  B   s  B    �    �   s  B   s      B  , ,  B  �  B  �  �  �  �  �  B  �      B  , ,  B  C  B  �  �  �  �  C  B  C      B  , ,  B  �  B  U  �  U  �  �  B  �      B  , ,  B    B  �  �  �  �    B        B  , ,  E  
K  E  
�  �  
�  �  
K  E  
K      B  , ,  E  �  E  ]  �  ]  �  �  E  �      B  , ,  E    E  �  �  �  �    E        B  , ,  E  �  E  -  �  -  �  �  E  �      B  , ,  E  �  E  �  �  �  �  �  E  �      B  , ,  E  S  E  �  �  �  �  S  E  S      B  , ,  E  �  E  e  �  e  �  �  E  �      B  , ,  B  {  B  %  �  %  �  {  B  {      B  , ,  B  �  B  	�  �  	�  �  �  B  �      B  , ,  B  
K  B  
�  �  
�  �  
K  B  
K      B  , ,  B  �  B  ]  �  ]  �  �  B  �      B  , ,  B    B  �  �  �  �    B        B  , ,  B  �  B  -  �  -  �  �  B  �      B  , ,  B  �  B  �  �  �  �  �  B  �      B  , ,  B  S  B  �  �  �  �  S  B  S      B  , ,  B  �  B  e  �  e  �  �  B  �      B  , ,  r  �  r  U    U    �  r  �      B  , ,  r    r  �    �      r        B  , ,  r  {  r  %    %    {  r  {      B  , ,  r  �  r  	�    	�    �  r  �      B  , ,  r  
K  r  
�    
�    
K  r  
K      B  , ,  r  �  r  ]    ]    �  r  �      B  , ,  r    r  �    �      r        B  , ,  r  �  r  -    -    �  r  �      B  , ,  r  �  r  �    �    �  r  �      B  , ,  r  S  r  �    �    S  r  S      B  , ,  r  �  r  e    e    �  r  �      B  , ,  �   s  �    W    W   s  �   s      B  , ,  �  �  �  �  W  �  W  �  �  �      B  , ,  r   s  r           s  r   s      B  , ,  �  C  �  �  W  �  W  C  �  C      B  , ,  �  �  �  U  W  U  W  �  �  �      B  , ,  �    �  �  W  �  W    �        B  , ,  �  {  �  %  W  %  W  {  �  {      B  , ,  �  �  �  	�  W  	�  W  �  �  �      B  , ,  �  
K  �  
�  W  
�  W  
K  �  
K      B  , ,  �  �  �  ]  W  ]  W  �  �  �      B  , ,  �    �  �  W  �  W    �        B  , ,  �  �  �  -  W  -  W  �  �  �      B  , ,  �  �  �  �  W  �  W  �  �  �      B  , ,  �  S  �  �  W  �  W  S  �  S      B  , ,  �  �  �  e  W  e  W  �  �  �      B  , ,  r  �  r  �    �    �  r  �      B  , ,  r  C  r  �    �    C  r  C      B  , ,  E   s  E    �    �   s  E   s      B  , ,  E  �  E  �  �  �  �  �  E  �      B  , ,  E  C  E  �  �  �  �  C  E  C      B  , ,  E  �  E  U  �  U  �  �  E  �      B  , ,  E    E  �  �  �  �    E        B  , ,  E  {  E  %  �  %  �  {  E  {      B  , ,  �   s  �    �    �   s  �   s      B  , ,  �  �  �  �  �  �  �  �  �  �      B  , ,  �  C  �  �  �  �  �  C  �  C      B  , ,  �  �  �  U  �  U  �  �  �  �      B  , ,  �    �  �  �  �  �    �        A   ,              �@  �  �@  �                  ]  , ,  �����  �  ��  D  ��  D����  �����      @   ,������������  �  �  �  �������������     � 
   % 0� 
   % 0 nfet$10     B   ,  ����8  �  u�  
d  u�  
d���8  ����8      B   ,  �  u�  �  wB  
d  wB  
d  u�  �  u�      D   ,   #   _   #  t�  q  t�  q   _   #   _      D   ,  
�   _  
�  t�  �  t�  �   _  
�   _      D   ,    v*    w  	�  w  	�  v*    v*      _   ,  �  u�  �  wL  
n  wL  
n  u�  �  u�      C   ,   A   K   A  t�  S  t�  S   K   A   K      C   ,  
�   K  
�  t�  �  t�  �   K  
�   K      C   ,    vH    v�  	�  v�  	�  vH    vH      C  , ,   A  ;�   A  <U   �  <U   �  ;�   A  ;�      C  , ,  �  ;�  �  <U  S  <U  S  ;�  �  ;�      C  , ,  
�  ;�  
�  <U  O  <U  O  ;�  
�  ;�      C  , ,    ;�    <U  �  <U  �  ;�    ;�      C  , ,   A  Y3   A  Y�   �  Y�   �  Y3   A  Y3      C  , ,  �  Y3  �  Y�  S  Y�  S  Y3  �  Y3      C  , ,  
�  Y3  
�  Y�  O  Y�  O  Y3  
�  Y3      C  , ,    Y3    Y�  �  Y�  �  Y3    Y3      C  , ,   A  ^�   A  _}   �  _}   �  ^�   A  ^�      C  , ,   A  `;   A  `�   �  `�   �  `;   A  `;      C  , ,   A  a�   A  bM   �  bM   �  a�   A  a�      C  , ,   A  c   A  c�   �  c�   �  c   A  c      C  , ,   A  ds   A  e   �  e   �  ds   A  ds      C  , ,   A  e�   A  f�   �  f�   �  e�   A  e�      C  , ,   A  gC   A  g�   �  g�   �  gC   A  gC      C  , ,   A  h�   A  iU   �  iU   �  h�   A  h�      C  , ,   A  j   A  j�   �  j�   �  j   A  j      C  , ,   A  k{   A  l%   �  l%   �  k{   A  k{      C  , ,   A  l�   A  m�   �  m�   �  l�   A  l�      C  , ,   A  nK   A  n�   �  n�   �  nK   A  nK      C  , ,   A  o�   A  p]   �  p]   �  o�   A  o�      C  , ,   A  q   A  q�   �  q�   �  q   A  q      C  , ,   A  r�   A  s-   �  s-   �  r�   A  r�      C  , ,   A  s�   A  t�   �  t�   �  s�   A  s�      C  , ,   A  Z�   A  [E   �  [E   �  Z�   A  Z�      C  , ,  �  Z�  �  [E  S  [E  S  Z�  �  Z�      C  , ,  �  \  �  \�  S  \�  S  \  �  \      C  , ,  �  ]k  �  ^  S  ^  S  ]k  �  ]k      C  , ,  �  ^�  �  _}  S  _}  S  ^�  �  ^�      C  , ,  �  `;  �  `�  S  `�  S  `;  �  `;      C  , ,  �  a�  �  bM  S  bM  S  a�  �  a�      C  , ,  �  c  �  c�  S  c�  S  c  �  c      C  , ,  �  ds  �  e  S  e  S  ds  �  ds      C  , ,  �  e�  �  f�  S  f�  S  e�  �  e�      C  , ,  �  gC  �  g�  S  g�  S  gC  �  gC      C  , ,  �  h�  �  iU  S  iU  S  h�  �  h�      C  , ,  �  j  �  j�  S  j�  S  j  �  j      C  , ,  �  k{  �  l%  S  l%  S  k{  �  k{      C  , ,  �  l�  �  m�  S  m�  S  l�  �  l�      C  , ,  �  nK  �  n�  S  n�  S  nK  �  nK      C  , ,  �  o�  �  p]  S  p]  S  o�  �  o�      C  , ,  �  q  �  q�  S  q�  S  q  �  q      C  , ,  �  r�  �  s-  S  s-  S  r�  �  r�      C  , ,  �  s�  �  t�  S  t�  S  s�  �  s�      C  , ,   A  \   A  \�   �  \�   �  \   A  \      C  , ,  
�  Z�  
�  [E  O  [E  O  Z�  
�  Z�      C  , ,  
�  \  
�  \�  O  \�  O  \  
�  \      C  , ,  
�  ]k  
�  ^  O  ^  O  ]k  
�  ]k      C  , ,  
�  ^�  
�  _}  O  _}  O  ^�  
�  ^�      C  , ,  
�  `;  
�  `�  O  `�  O  `;  
�  `;      C  , ,  
�  a�  
�  bM  O  bM  O  a�  
�  a�      C  , ,  
�  c  
�  c�  O  c�  O  c  
�  c      C  , ,  
�  ds  
�  e  O  e  O  ds  
�  ds      C  , ,  
�  e�  
�  f�  O  f�  O  e�  
�  e�      C  , ,  
�  gC  
�  g�  O  g�  O  gC  
�  gC      C  , ,  
�  h�  
�  iU  O  iU  O  h�  
�  h�      C  , ,  
�  j  
�  j�  O  j�  O  j  
�  j      C  , ,  
�  k{  
�  l%  O  l%  O  k{  
�  k{      C  , ,  
�  l�  
�  m�  O  m�  O  l�  
�  l�      C  , ,  
�  nK  
�  n�  O  n�  O  nK  
�  nK      C  , ,  
�  o�  
�  p]  O  p]  O  o�  
�  o�      C  , ,  
�  q  
�  q�  O  q�  O  q  
�  q      C  , ,  
�  r�  
�  s-  O  s-  O  r�  
�  r�      C  , ,  
�  s�  
�  t�  O  t�  O  s�  
�  s�      C  , ,   A  ]k   A  ^   �  ^   �  ]k   A  ]k      C  , ,    Z�    [E  �  [E  �  Z�    Z�      C  , ,    \    \�  �  \�  �  \    \      C  , ,    ]k    ^  �  ^  �  ]k    ]k      C  , ,    ^�    _}  �  _}  �  ^�    ^�      C  , ,    `;    `�  �  `�  �  `;    `;      C  , ,    a�    bM  �  bM  �  a�    a�      C  , ,    c    c�  �  c�  �  c    c      C  , ,    ds    e  �  e  �  ds    ds      C  , ,    e�    f�  �  f�  �  e�    e�      C  , ,    gC    g�  �  g�  �  gC    gC      C  , ,    h�    iU  �  iU  �  h�    h�      C  , ,    j    j�  �  j�  �  j    j      C  , ,    k{    l%  �  l%  �  k{    k{      C  , ,    l�    m�  �  m�  �  l�    l�      C  , ,    nK    n�  �  n�  �  nK    nK      C  , ,    o�    p]  �  p]  �  o�    o�      C  , ,    q    q�  �  q�  �  q    q      C  , ,    r�    s-  �  s-  �  r�    r�      C  , ,    s�    t�  �  t�  �  s�    s�      C  , ,  W  vH  W  v�    v�    vH  W  vH      C  , ,  �  vH  �  v�  i  v�  i  vH  �  vH      C  , ,  '  vH  '  v�  �  v�  �  vH  '  vH      C  , ,  �  vH  �  v�  9  v�  9  vH  �  vH      C  , ,  �  vH  �  v�  	�  v�  	�  vH  �  vH      C  , ,  
�  E�  
�  F-  O  F-  O  E�  
�  E�      C  , ,  
�  F�  
�  G�  O  G�  O  F�  
�  F�      C  , ,  
�  HS  
�  H�  O  H�  O  HS  
�  HS      C  , ,  
�  I�  
�  Je  O  Je  O  I�  
�  I�      C  , ,  
�  K#  
�  K�  O  K�  O  K#  
�  K#      C  , ,  
�  L�  
�  M5  O  M5  O  L�  
�  L�      C  , ,  
�  M�  
�  N�  O  N�  O  M�  
�  M�      C  , ,  
�  O[  
�  P  O  P  O  O[  
�  O[      C  , ,  
�  P�  
�  Qm  O  Qm  O  P�  
�  P�      C  , ,  
�  R+  
�  R�  O  R�  O  R+  
�  R+      C  , ,  
�  S�  
�  T=  O  T=  O  S�  
�  S�      C  , ,  
�  T�  
�  U�  O  U�  O  T�  
�  T�      C  , ,  
�  Vc  
�  W  O  W  O  Vc  
�  Vc      C  , ,  
�  W�  
�  Xu  O  Xu  O  W�  
�  W�      C  , ,  �  ?�  �  @�  S  @�  S  ?�  �  ?�      C  , ,  �  AK  �  A�  S  A�  S  AK  �  AK      C  , ,  �  B�  �  C]  S  C]  S  B�  �  B�      C  , ,  �  D  �  D�  S  D�  S  D  �  D      C  , ,  �  E�  �  F-  S  F-  S  E�  �  E�      C  , ,  �  F�  �  G�  S  G�  S  F�  �  F�      C  , ,  �  HS  �  H�  S  H�  S  HS  �  HS      C  , ,  �  I�  �  Je  S  Je  S  I�  �  I�      C  , ,  �  K#  �  K�  S  K�  S  K#  �  K#      C  , ,  �  L�  �  M5  S  M5  S  L�  �  L�      C  , ,  �  M�  �  N�  S  N�  S  M�  �  M�      C  , ,  �  O[  �  P  S  P  S  O[  �  O[      C  , ,  �  P�  �  Qm  S  Qm  S  P�  �  P�      C  , ,  �  R+  �  R�  S  R�  S  R+  �  R+      C  , ,  �  S�  �  T=  S  T=  S  S�  �  S�      C  , ,  �  T�  �  U�  S  U�  S  T�  �  T�      C  , ,  �  Vc  �  W  S  W  S  Vc  �  Vc      C  , ,  �  W�  �  Xu  S  Xu  S  W�  �  W�      C  , ,   A  E�   A  F-   �  F-   �  E�   A  E�      C  , ,   A  F�   A  G�   �  G�   �  F�   A  F�      C  , ,   A  ?�   A  @�   �  @�   �  ?�   A  ?�      C  , ,    =    =�  �  =�  �  =    =      C  , ,    >{    ?%  �  ?%  �  >{    >{      C  , ,    ?�    @�  �  @�  �  ?�    ?�      C  , ,    AK    A�  �  A�  �  AK    AK      C  , ,    B�    C]  �  C]  �  B�    B�      C  , ,    D    D�  �  D�  �  D    D      C  , ,    E�    F-  �  F-  �  E�    E�      C  , ,    F�    G�  �  G�  �  F�    F�      C  , ,    HS    H�  �  H�  �  HS    HS      C  , ,    I�    Je  �  Je  �  I�    I�      C  , ,    K#    K�  �  K�  �  K#    K#      C  , ,    L�    M5  �  M5  �  L�    L�      C  , ,    M�    N�  �  N�  �  M�    M�      C  , ,    O[    P  �  P  �  O[    O[      C  , ,    P�    Qm  �  Qm  �  P�    P�      C  , ,    R+    R�  �  R�  �  R+    R+      C  , ,    S�    T=  �  T=  �  S�    S�      C  , ,    T�    U�  �  U�  �  T�    T�      C  , ,    Vc    W  �  W  �  Vc    Vc      C  , ,    W�    Xu  �  Xu  �  W�    W�      C  , ,   A  HS   A  H�   �  H�   �  HS   A  HS      C  , ,   A  I�   A  Je   �  Je   �  I�   A  I�      C  , ,   A  K#   A  K�   �  K�   �  K#   A  K#      C  , ,   A  L�   A  M5   �  M5   �  L�   A  L�      C  , ,   A  M�   A  N�   �  N�   �  M�   A  M�      C  , ,   A  O[   A  P   �  P   �  O[   A  O[      C  , ,   A  P�   A  Qm   �  Qm   �  P�   A  P�      C  , ,   A  R+   A  R�   �  R�   �  R+   A  R+      C  , ,   A  S�   A  T=   �  T=   �  S�   A  S�      C  , ,   A  T�   A  U�   �  U�   �  T�   A  T�      C  , ,   A  Vc   A  W   �  W   �  Vc   A  Vc      C  , ,   A  W�   A  Xu   �  Xu   �  W�   A  W�      C  , ,   A  AK   A  A�   �  A�   �  AK   A  AK      C  , ,   A  B�   A  C]   �  C]   �  B�   A  B�      C  , ,   A  D   A  D�   �  D�   �  D   A  D      C  , ,   A  =   A  =�   �  =�   �  =   A  =      C  , ,  �  =  �  =�  S  =�  S  =  �  =      C  , ,  �  >{  �  ?%  S  ?%  S  >{  �  >{      C  , ,   A  >{   A  ?%   �  ?%   �  >{   A  >{      C  , ,  
�  =  
�  =�  O  =�  O  =  
�  =      C  , ,  
�  >{  
�  ?%  O  ?%  O  >{  
�  >{      C  , ,  
�  ?�  
�  @�  O  @�  O  ?�  
�  ?�      C  , ,  
�  AK  
�  A�  O  A�  O  AK  
�  AK      C  , ,  
�  B�  
�  C]  O  C]  O  B�  
�  B�      C  , ,  
�  D  
�  D�  O  D�  O  D  
�  D      C  , ,  
�  #  
�  �  O  �  O  #  
�  #      C  , ,  �  #  �  �  S  �  S  #  �  #      C  , ,    #    �  �  �  �  #    #      C  , ,   A  #   A  �   �  �   �  #   A  #      C  , ,  
�  #�  
�  $m  O  $m  O  #�  
�  #�      C  , ,  
�  %+  
�  %�  O  %�  O  %+  
�  %+      C  , ,  
�  &�  
�  '=  O  '=  O  &�  
�  &�      C  , ,  
�  '�  
�  (�  O  (�  O  '�  
�  '�      C  , ,  
�  )c  
�  *  O  *  O  )c  
�  )c      C  , ,  
�  *�  
�  +u  O  +u  O  *�  
�  *�      C  , ,  
�  ,3  
�  ,�  O  ,�  O  ,3  
�  ,3      C  , ,  
�  -�  
�  .E  O  .E  O  -�  
�  -�      C  , ,  
�  /  
�  /�  O  /�  O  /  
�  /      C  , ,  
�  0k  
�  1  O  1  O  0k  
�  0k      C  , ,  
�  1�  
�  2}  O  2}  O  1�  
�  1�      C  , ,  
�  3;  
�  3�  O  3�  O  3;  
�  3;      C  , ,  
�  4�  
�  5M  O  5M  O  4�  
�  4�      C  , ,  
�  6  
�  6�  O  6�  O  6  
�  6      C  , ,  
�  7s  
�  8  O  8  O  7s  
�  7s      C  , ,  
�  8�  
�  9�  O  9�  O  8�  
�  8�      C  , ,  
�  :C  
�  :�  O  :�  O  :C  
�  :C      C  , ,   A  8�   A  9�   �  9�   �  8�   A  8�      C  , ,  
�  �  
�   5  O   5  O  �  
�  �      C  , ,  �  �  �   5  S   5  S  �  �  �      C  , ,  �   �  �  !�  S  !�  S   �  �   �      C  , ,  �  "[  �  #  S  #  S  "[  �  "[      C  , ,  �  #�  �  $m  S  $m  S  #�  �  #�      C  , ,  �  %+  �  %�  S  %�  S  %+  �  %+      C  , ,  �  &�  �  '=  S  '=  S  &�  �  &�      C  , ,  �  '�  �  (�  S  (�  S  '�  �  '�      C  , ,  �  )c  �  *  S  *  S  )c  �  )c      C  , ,  �  *�  �  +u  S  +u  S  *�  �  *�      C  , ,  �  ,3  �  ,�  S  ,�  S  ,3  �  ,3      C  , ,  �  -�  �  .E  S  .E  S  -�  �  -�      C  , ,  �  /  �  /�  S  /�  S  /  �  /      C  , ,  �  0k  �  1  S  1  S  0k  �  0k      C  , ,  �  1�  �  2}  S  2}  S  1�  �  1�      C  , ,  �  3;  �  3�  S  3�  S  3;  �  3;      C  , ,  �  4�  �  5M  S  5M  S  4�  �  4�      C  , ,  �  6  �  6�  S  6�  S  6  �  6      C  , ,  �  7s  �  8  S  8  S  7s  �  7s      C  , ,  
�   �  
�  !�  O  !�  O   �  
�   �      C  , ,    �     5  �   5  �  �    �      C  , ,     �    !�  �  !�  �   �     �      C  , ,    "[    #  �  #  �  "[    "[      C  , ,    #�    $m  �  $m  �  #�    #�      C  , ,    %+    %�  �  %�  �  %+    %+      C  , ,    &�    '=  �  '=  �  &�    &�      C  , ,    '�    (�  �  (�  �  '�    '�      C  , ,    )c    *  �  *  �  )c    )c      C  , ,    *�    +u  �  +u  �  *�    *�      C  , ,    ,3    ,�  �  ,�  �  ,3    ,3      C  , ,    -�    .E  �  .E  �  -�    -�      C  , ,    /    /�  �  /�  �  /    /      C  , ,    0k    1  �  1  �  0k    0k      C  , ,    1�    2}  �  2}  �  1�    1�      C  , ,    3;    3�  �  3�  �  3;    3;      C  , ,    4�    5M  �  5M  �  4�    4�      C  , ,    6    6�  �  6�  �  6    6      C  , ,    7s    8  �  8  �  7s    7s      C  , ,    8�    9�  �  9�  �  8�    8�      C  , ,    :C    :�  �  :�  �  :C    :C      C  , ,  �  8�  �  9�  S  9�  S  8�  �  8�      C  , ,  �  :C  �  :�  S  :�  S  :C  �  :C      C  , ,   A  :C   A  :�   �  :�   �  :C   A  :C      C  , ,  
�  "[  
�  #  O  #  O  "[  
�  "[      C  , ,   A  �   A   5   �   5   �  �   A  �      C  , ,   A   �   A  !�   �  !�   �   �   A   �      C  , ,   A  "[   A  #   �  #   �  "[   A  "[      C  , ,   A  #�   A  $m   �  $m   �  #�   A  #�      C  , ,   A  %+   A  %�   �  %�   �  %+   A  %+      C  , ,   A  &�   A  '=   �  '=   �  &�   A  &�      C  , ,   A  '�   A  (�   �  (�   �  '�   A  '�      C  , ,   A  )c   A  *   �  *   �  )c   A  )c      C  , ,   A  *�   A  +u   �  +u   �  *�   A  *�      C  , ,   A  ,3   A  ,�   �  ,�   �  ,3   A  ,3      C  , ,   A  -�   A  .E   �  .E   �  -�   A  -�      C  , ,   A  /   A  /�   �  /�   �  /   A  /      C  , ,   A  0k   A  1   �  1   �  0k   A  0k      C  , ,   A  1�   A  2}   �  2}   �  1�   A  1�      C  , ,   A  3;   A  3�   �  3�   �  3;   A  3;      C  , ,   A  4�   A  5M   �  5M   �  4�   A  4�      C  , ,   A  6   A  6�   �  6�   �  6   A  6      C  , ,   A  7s   A  8   �  8   �  7s   A  7s      C  , ,    ;    �  �  �  �  ;    ;      C  , ,    �    M  �  M  �  �    �      C  , ,    	    	�  �  	�  �  	    	      C  , ,    
s      �    �  
s    
s      C  , ,    �    �  �  �  �  �    �      C  , ,    C    �  �  �  �  C    C      C  , ,    �    U  �  U  �  �    �      C  , ,        �  �  �  �            C  , ,    {    %  �  %  �  {    {      C  , ,    �    �  �  �  �  �    �      C  , ,    K    �  �  �  �  K    K      C  , ,    �    ]  �  ]  �  �    �      C  , ,        �  �  �  �            C  , ,    �    -  �  -  �  �    �      C  , ,    �    �  �  �  �  �    �      C  , ,    S    �  �  �  �  S    S      C  , ,    �    e  �  e  �  �    �      C  , ,  �    �  �  S  �  S    �        C  , ,  �  k  �    S    S  k  �  k      C  , ,  �  �  �  }  S  }  S  �  �  �      C  , ,  �  ;  �  �  S  �  S  ;  �  ;      C  , ,  �  �  �  M  S  M  S  �  �  �      C  , ,  �  	  �  	�  S  	�  S  	  �  	      C  , ,  �  
s  �    S    S  
s  �  
s      C  , ,  �  �  �  �  S  �  S  �  �  �      C  , ,  �  C  �  �  S  �  S  C  �  C      C  , ,  �  �  �  U  S  U  S  �  �  �      C  , ,  �    �  �  S  �  S    �        C  , ,  �  {  �  %  S  %  S  {  �  {      C  , ,  �  �  �  �  S  �  S  �  �  �      C  , ,  �  K  �  �  S  �  S  K  �  K      C  , ,  �  �  �  ]  S  ]  S  �  �  �      C  , ,  �    �  �  S  �  S    �        C  , ,  �  �  �  -  S  -  S  �  �  �      C  , ,  �  �  �  �  S  �  S  �  �  �      C  , ,  �  S  �  �  S  �  S  S  �  S      C  , ,  �  �  �  e  S  e  S  �  �  �      C  , ,  
�  
s  
�    O    O  
s  
�  
s      C  , ,  
�  �  
�  �  O  �  O  �  
�  �      C  , ,  
�  C  
�  �  O  �  O  C  
�  C      C  , ,  
�  �  
�  U  O  U  O  �  
�  �      C  , ,   A   �   A  E   �  E   �   �   A   �      C  , ,   A     A  �   �  �   �     A        C  , ,   A  k   A     �     �  k   A  k      C  , ,   A  �   A  }   �  }   �  �   A  �      C  , ,   A  ;   A  �   �  �   �  ;   A  ;      C  , ,   A  �   A  M   �  M   �  �   A  �      C  , ,   A  	   A  	�   �  	�   �  	   A  	      C  , ,   A  
s   A     �     �  
s   A  
s      C  , ,   A  �   A  �   �  �   �  �   A  �      C  , ,   A  C   A  �   �  �   �  C   A  C      C  , ,   A  �   A  U   �  U   �  �   A  �      C  , ,   A     A  �   �  �   �     A        C  , ,   A  {   A  %   �  %   �  {   A  {      C  , ,   A  �   A  �   �  �   �  �   A  �      C  , ,   A  K   A  �   �  �   �  K   A  K      C  , ,   A  �   A  ]   �  ]   �  �   A  �      C  , ,   A     A  �   �  �   �     A        C  , ,   A  �   A  -   �  -   �  �   A  �      C  , ,   A  �   A  �   �  �   �  �   A  �      C  , ,   A  S   A  �   �  �   �  S   A  S      C  , ,   A  �   A  e   �  e   �  �   A  �      C  , ,  
�    
�  �  O  �  O    
�        C  , ,  
�  {  
�  %  O  %  O  {  
�  {      C  , ,  
�  �  
�  �  O  �  O  �  
�  �      C  , ,  
�  K  
�  �  O  �  O  K  
�  K      C  , ,  
�  �  
�  ]  O  ]  O  �  
�  �      C  , ,  
�    
�  �  O  �  O    
�        C  , ,  
�  �  
�  -  O  -  O  �  
�  �      C  , ,  
�  �  
�  �  O  �  O  �  
�  �      C  , ,  
�  S  
�  �  O  �  O  S  
�  S      C  , ,  
�  �  
�  e  O  e  O  �  
�  �      C  , ,  
�  �  
�  }  O  }  O  �  
�  �      C  , ,  
�  ;  
�  �  O  �  O  ;  
�  ;      C  , ,  
�  �  
�  M  O  M  O  �  
�  �      C  , ,  
�  	  
�  	�  O  	�  O  	  
�  	      C  , ,  �   �  �  E  S  E  S   �  �   �      C  , ,     �    E  �  E  �   �     �      C  , ,        �  �  �  �            C  , ,    k      �    �  k    k      C  , ,    �    }  �  }  �  �    �      C  , ,  
�   �  
�  E  O  E  O   �  
�   �      C  , ,  
�    
�  �  O  �  O    
�        C  , ,  
�  k  
�    O    O  k  
�  k      B  , ,   A  ;�   A  <U   �  <U   �  ;�   A  ;�      B  , ,  �  ;�  �  <U  S  <U  S  ;�  �  ;�      B  , ,  
�  ;�  
�  <U  O  <U  O  ;�  
�  ;�      B  , ,    ;�    <U  �  <U  �  ;�    ;�      B  , ,   A  Y3   A  Y�   �  Y�   �  Y3   A  Y3      B  , ,  �  Y3  �  Y�  S  Y�  S  Y3  �  Y3      B  , ,  
�  Y3  
�  Y�  O  Y�  O  Y3  
�  Y3      B  , ,    Y3    Y�  �  Y�  �  Y3    Y3      B  , ,   A  ^�   A  _}   �  _}   �  ^�   A  ^�      B  , ,   A  `;   A  `�   �  `�   �  `;   A  `;      B  , ,   A  a�   A  bM   �  bM   �  a�   A  a�      B  , ,   A  c   A  c�   �  c�   �  c   A  c      B  , ,   A  ds   A  e   �  e   �  ds   A  ds      B  , ,   A  e�   A  f�   �  f�   �  e�   A  e�      B  , ,   A  gC   A  g�   �  g�   �  gC   A  gC      B  , ,   A  h�   A  iU   �  iU   �  h�   A  h�      B  , ,   A  j   A  j�   �  j�   �  j   A  j      B  , ,   A  k{   A  l%   �  l%   �  k{   A  k{      B  , ,   A  l�   A  m�   �  m�   �  l�   A  l�      B  , ,   A  nK   A  n�   �  n�   �  nK   A  nK      B  , ,   A  o�   A  p]   �  p]   �  o�   A  o�      B  , ,   A  q   A  q�   �  q�   �  q   A  q      B  , ,   A  r�   A  s-   �  s-   �  r�   A  r�      B  , ,   A  s�   A  t�   �  t�   �  s�   A  s�      B  , ,   A  Z�   A  [E   �  [E   �  Z�   A  Z�      B  , ,  �  Z�  �  [E  S  [E  S  Z�  �  Z�      B  , ,  �  \  �  \�  S  \�  S  \  �  \      B  , ,  �  ]k  �  ^  S  ^  S  ]k  �  ]k      B  , ,  �  ^�  �  _}  S  _}  S  ^�  �  ^�      B  , ,  �  `;  �  `�  S  `�  S  `;  �  `;      B  , ,  �  a�  �  bM  S  bM  S  a�  �  a�      B  , ,  �  c  �  c�  S  c�  S  c  �  c      B  , ,  �  ds  �  e  S  e  S  ds  �  ds      B  , ,  �  e�  �  f�  S  f�  S  e�  �  e�      B  , ,  �  gC  �  g�  S  g�  S  gC  �  gC      B  , ,  �  h�  �  iU  S  iU  S  h�  �  h�      B  , ,  �  j  �  j�  S  j�  S  j  �  j      B  , ,  �  k{  �  l%  S  l%  S  k{  �  k{      B  , ,  �  l�  �  m�  S  m�  S  l�  �  l�      B  , ,  �  nK  �  n�  S  n�  S  nK  �  nK      B  , ,  �  o�  �  p]  S  p]  S  o�  �  o�      B  , ,  �  q  �  q�  S  q�  S  q  �  q      B  , ,  �  r�  �  s-  S  s-  S  r�  �  r�      B  , ,  �  s�  �  t�  S  t�  S  s�  �  s�      B  , ,   A  \   A  \�   �  \�   �  \   A  \      B  , ,  
�  Z�  
�  [E  O  [E  O  Z�  
�  Z�      B  , ,  
�  \  
�  \�  O  \�  O  \  
�  \      B  , ,  
�  ]k  
�  ^  O  ^  O  ]k  
�  ]k      B  , ,  
�  ^�  
�  _}  O  _}  O  ^�  
�  ^�      B  , ,  
�  `;  
�  `�  O  `�  O  `;  
�  `;      B  , ,  
�  a�  
�  bM  O  bM  O  a�  
�  a�      B  , ,  
�  c  
�  c�  O  c�  O  c  
�  c      B  , ,  
�  ds  
�  e  O  e  O  ds  
�  ds      B  , ,  
�  e�  
�  f�  O  f�  O  e�  
�  e�      B  , ,  
�  gC  
�  g�  O  g�  O  gC  
�  gC      B  , ,  
�  h�  
�  iU  O  iU  O  h�  
�  h�      B  , ,  
�  j  
�  j�  O  j�  O  j  
�  j      B  , ,  
�  k{  
�  l%  O  l%  O  k{  
�  k{      B  , ,  
�  l�  
�  m�  O  m�  O  l�  
�  l�      B  , ,  
�  nK  
�  n�  O  n�  O  nK  
�  nK      B  , ,  
�  o�  
�  p]  O  p]  O  o�  
�  o�      B  , ,  
�  q  
�  q�  O  q�  O  q  
�  q      B  , ,  
�  r�  
�  s-  O  s-  O  r�  
�  r�      B  , ,  
�  s�  
�  t�  O  t�  O  s�  
�  s�      B  , ,   A  ]k   A  ^   �  ^   �  ]k   A  ]k      B  , ,    Z�    [E  �  [E  �  Z�    Z�      B  , ,    \    \�  �  \�  �  \    \      B  , ,    ]k    ^  �  ^  �  ]k    ]k      B  , ,    ^�    _}  �  _}  �  ^�    ^�      B  , ,    `;    `�  �  `�  �  `;    `;      B  , ,    a�    bM  �  bM  �  a�    a�      B  , ,    c    c�  �  c�  �  c    c      B  , ,    ds    e  �  e  �  ds    ds      B  , ,    e�    f�  �  f�  �  e�    e�      B  , ,    gC    g�  �  g�  �  gC    gC      B  , ,    h�    iU  �  iU  �  h�    h�      B  , ,    j    j�  �  j�  �  j    j      B  , ,    k{    l%  �  l%  �  k{    k{      B  , ,    l�    m�  �  m�  �  l�    l�      B  , ,    nK    n�  �  n�  �  nK    nK      B  , ,    o�    p]  �  p]  �  o�    o�      B  , ,    q    q�  �  q�  �  q    q      B  , ,    r�    s-  �  s-  �  r�    r�      B  , ,    s�    t�  �  t�  �  s�    s�      B  , ,  W  vH  W  v�    v�    vH  W  vH      B  , ,  �  vH  �  v�  i  v�  i  vH  �  vH      B  , ,  '  vH  '  v�  �  v�  �  vH  '  vH      B  , ,  �  vH  �  v�  9  v�  9  vH  �  vH      B  , ,  �  vH  �  v�  	�  v�  	�  vH  �  vH      B  , ,  
�  E�  
�  F-  O  F-  O  E�  
�  E�      B  , ,  
�  F�  
�  G�  O  G�  O  F�  
�  F�      B  , ,  
�  HS  
�  H�  O  H�  O  HS  
�  HS      B  , ,  
�  I�  
�  Je  O  Je  O  I�  
�  I�      B  , ,  
�  K#  
�  K�  O  K�  O  K#  
�  K#      B  , ,  
�  L�  
�  M5  O  M5  O  L�  
�  L�      B  , ,  
�  M�  
�  N�  O  N�  O  M�  
�  M�      B  , ,  
�  O[  
�  P  O  P  O  O[  
�  O[      B  , ,  
�  P�  
�  Qm  O  Qm  O  P�  
�  P�      B  , ,  
�  R+  
�  R�  O  R�  O  R+  
�  R+      B  , ,  
�  S�  
�  T=  O  T=  O  S�  
�  S�      B  , ,  
�  T�  
�  U�  O  U�  O  T�  
�  T�      B  , ,  
�  Vc  
�  W  O  W  O  Vc  
�  Vc      B  , ,  
�  W�  
�  Xu  O  Xu  O  W�  
�  W�      B  , ,  �  ?�  �  @�  S  @�  S  ?�  �  ?�      B  , ,  �  AK  �  A�  S  A�  S  AK  �  AK      B  , ,  �  B�  �  C]  S  C]  S  B�  �  B�      B  , ,  �  D  �  D�  S  D�  S  D  �  D      B  , ,  �  E�  �  F-  S  F-  S  E�  �  E�      B  , ,  �  F�  �  G�  S  G�  S  F�  �  F�      B  , ,  �  HS  �  H�  S  H�  S  HS  �  HS      B  , ,  �  I�  �  Je  S  Je  S  I�  �  I�      B  , ,  �  K#  �  K�  S  K�  S  K#  �  K#      B  , ,  �  L�  �  M5  S  M5  S  L�  �  L�      B  , ,  �  M�  �  N�  S  N�  S  M�  �  M�      B  , ,  �  O[  �  P  S  P  S  O[  �  O[      B  , ,  �  P�  �  Qm  S  Qm  S  P�  �  P�      B  , ,  �  R+  �  R�  S  R�  S  R+  �  R+      B  , ,  �  S�  �  T=  S  T=  S  S�  �  S�      B  , ,  �  T�  �  U�  S  U�  S  T�  �  T�      B  , ,  �  Vc  �  W  S  W  S  Vc  �  Vc      B  , ,  �  W�  �  Xu  S  Xu  S  W�  �  W�      B  , ,   A  E�   A  F-   �  F-   �  E�   A  E�      B  , ,   A  F�   A  G�   �  G�   �  F�   A  F�      B  , ,   A  ?�   A  @�   �  @�   �  ?�   A  ?�      B  , ,    =    =�  �  =�  �  =    =      B  , ,    >{    ?%  �  ?%  �  >{    >{      B  , ,    ?�    @�  �  @�  �  ?�    ?�      B  , ,    AK    A�  �  A�  �  AK    AK      B  , ,    B�    C]  �  C]  �  B�    B�      B  , ,    D    D�  �  D�  �  D    D      B  , ,    E�    F-  �  F-  �  E�    E�      B  , ,    F�    G�  �  G�  �  F�    F�      B  , ,    HS    H�  �  H�  �  HS    HS      B  , ,    I�    Je  �  Je  �  I�    I�      B  , ,    K#    K�  �  K�  �  K#    K#      B  , ,    L�    M5  �  M5  �  L�    L�      B  , ,    M�    N�  �  N�  �  M�    M�      B  , ,    O[    P  �  P  �  O[    O[      B  , ,    P�    Qm  �  Qm  �  P�    P�      B  , ,    R+    R�  �  R�  �  R+    R+      B  , ,    S�    T=  �  T=  �  S�    S�      B  , ,    T�    U�  �  U�  �  T�    T�      B  , ,    Vc    W  �  W  �  Vc    Vc      B  , ,    W�    Xu  �  Xu  �  W�    W�      B  , ,   A  HS   A  H�   �  H�   �  HS   A  HS      B  , ,   A  I�   A  Je   �  Je   �  I�   A  I�      B  , ,   A  K#   A  K�   �  K�   �  K#   A  K#      B  , ,   A  L�   A  M5   �  M5   �  L�   A  L�      B  , ,   A  M�   A  N�   �  N�   �  M�   A  M�      B  , ,   A  O[   A  P   �  P   �  O[   A  O[      B  , ,   A  P�   A  Qm   �  Qm   �  P�   A  P�      B  , ,   A  R+   A  R�   �  R�   �  R+   A  R+      B  , ,   A  S�   A  T=   �  T=   �  S�   A  S�      B  , ,   A  T�   A  U�   �  U�   �  T�   A  T�      B  , ,   A  Vc   A  W   �  W   �  Vc   A  Vc      B  , ,   A  W�   A  Xu   �  Xu   �  W�   A  W�      B  , ,   A  AK   A  A�   �  A�   �  AK   A  AK      B  , ,   A  B�   A  C]   �  C]   �  B�   A  B�      B  , ,   A  D   A  D�   �  D�   �  D   A  D      B  , ,   A  =   A  =�   �  =�   �  =   A  =      B  , ,  �  =  �  =�  S  =�  S  =  �  =      B  , ,  �  >{  �  ?%  S  ?%  S  >{  �  >{      B  , ,   A  >{   A  ?%   �  ?%   �  >{   A  >{      B  , ,  
�  =  
�  =�  O  =�  O  =  
�  =      B  , ,  
�  >{  
�  ?%  O  ?%  O  >{  
�  >{      B  , ,  
�  ?�  
�  @�  O  @�  O  ?�  
�  ?�      B  , ,  
�  AK  
�  A�  O  A�  O  AK  
�  AK      B  , ,  
�  B�  
�  C]  O  C]  O  B�  
�  B�      B  , ,  
�  D  
�  D�  O  D�  O  D  
�  D      B  , ,  
�  #  
�  �  O  �  O  #  
�  #      B  , ,  �  #  �  �  S  �  S  #  �  #      B  , ,    #    �  �  �  �  #    #      B  , ,   A  #   A  �   �  �   �  #   A  #      B  , ,  
�  #�  
�  $m  O  $m  O  #�  
�  #�      B  , ,  
�  %+  
�  %�  O  %�  O  %+  
�  %+      B  , ,  
�  &�  
�  '=  O  '=  O  &�  
�  &�      B  , ,  
�  '�  
�  (�  O  (�  O  '�  
�  '�      B  , ,  
�  )c  
�  *  O  *  O  )c  
�  )c      B  , ,  
�  *�  
�  +u  O  +u  O  *�  
�  *�      B  , ,  
�  ,3  
�  ,�  O  ,�  O  ,3  
�  ,3      B  , ,  
�  -�  
�  .E  O  .E  O  -�  
�  -�      B  , ,  
�  /  
�  /�  O  /�  O  /  
�  /      B  , ,  
�  0k  
�  1  O  1  O  0k  
�  0k      B  , ,  
�  1�  
�  2}  O  2}  O  1�  
�  1�      B  , ,  
�  3;  
�  3�  O  3�  O  3;  
�  3;      B  , ,  
�  4�  
�  5M  O  5M  O  4�  
�  4�      B  , ,  
�  6  
�  6�  O  6�  O  6  
�  6      B  , ,  
�  7s  
�  8  O  8  O  7s  
�  7s      B  , ,  
�  8�  
�  9�  O  9�  O  8�  
�  8�      B  , ,  
�  :C  
�  :�  O  :�  O  :C  
�  :C      B  , ,   A  8�   A  9�   �  9�   �  8�   A  8�      B  , ,  
�  �  
�   5  O   5  O  �  
�  �      B  , ,  �  �  �   5  S   5  S  �  �  �      B  , ,  �   �  �  !�  S  !�  S   �  �   �      B  , ,  �  "[  �  #  S  #  S  "[  �  "[      B  , ,  �  #�  �  $m  S  $m  S  #�  �  #�      B  , ,  �  %+  �  %�  S  %�  S  %+  �  %+      B  , ,  �  &�  �  '=  S  '=  S  &�  �  &�      B  , ,  �  '�  �  (�  S  (�  S  '�  �  '�      B  , ,  �  )c  �  *  S  *  S  )c  �  )c      B  , ,  �  *�  �  +u  S  +u  S  *�  �  *�      B  , ,  �  ,3  �  ,�  S  ,�  S  ,3  �  ,3      B  , ,  �  -�  �  .E  S  .E  S  -�  �  -�      B  , ,  �  /  �  /�  S  /�  S  /  �  /      B  , ,  �  0k  �  1  S  1  S  0k  �  0k      B  , ,  �  1�  �  2}  S  2}  S  1�  �  1�      B  , ,  �  3;  �  3�  S  3�  S  3;  �  3;      B  , ,  �  4�  �  5M  S  5M  S  4�  �  4�      B  , ,  �  6  �  6�  S  6�  S  6  �  6      B  , ,  �  7s  �  8  S  8  S  7s  �  7s      B  , ,  
�   �  
�  !�  O  !�  O   �  
�   �      B  , ,    �     5  �   5  �  �    �      B  , ,     �    !�  �  !�  �   �     �      B  , ,    "[    #  �  #  �  "[    "[      B  , ,    #�    $m  �  $m  �  #�    #�      B  , ,    %+    %�  �  %�  �  %+    %+      B  , ,    &�    '=  �  '=  �  &�    &�      B  , ,    '�    (�  �  (�  �  '�    '�      B  , ,    )c    *  �  *  �  )c    )c      B  , ,    *�    +u  �  +u  �  *�    *�      B  , ,    ,3    ,�  �  ,�  �  ,3    ,3      B  , ,    -�    .E  �  .E  �  -�    -�      B  , ,    /    /�  �  /�  �  /    /      B  , ,    0k    1  �  1  �  0k    0k      B  , ,    1�    2}  �  2}  �  1�    1�      B  , ,    3;    3�  �  3�  �  3;    3;      B  , ,    4�    5M  �  5M  �  4�    4�      B  , ,    6    6�  �  6�  �  6    6      B  , ,    7s    8  �  8  �  7s    7s      B  , ,    8�    9�  �  9�  �  8�    8�      B  , ,    :C    :�  �  :�  �  :C    :C      B  , ,  �  8�  �  9�  S  9�  S  8�  �  8�      B  , ,  �  :C  �  :�  S  :�  S  :C  �  :C      B  , ,   A  :C   A  :�   �  :�   �  :C   A  :C      B  , ,  
�  "[  
�  #  O  #  O  "[  
�  "[      B  , ,   A  �   A   5   �   5   �  �   A  �      B  , ,   A   �   A  !�   �  !�   �   �   A   �      B  , ,   A  "[   A  #   �  #   �  "[   A  "[      B  , ,   A  #�   A  $m   �  $m   �  #�   A  #�      B  , ,   A  %+   A  %�   �  %�   �  %+   A  %+      B  , ,   A  &�   A  '=   �  '=   �  &�   A  &�      B  , ,   A  '�   A  (�   �  (�   �  '�   A  '�      B  , ,   A  )c   A  *   �  *   �  )c   A  )c      B  , ,   A  *�   A  +u   �  +u   �  *�   A  *�      B  , ,   A  ,3   A  ,�   �  ,�   �  ,3   A  ,3      B  , ,   A  -�   A  .E   �  .E   �  -�   A  -�      B  , ,   A  /   A  /�   �  /�   �  /   A  /      B  , ,   A  0k   A  1   �  1   �  0k   A  0k      B  , ,   A  1�   A  2}   �  2}   �  1�   A  1�      B  , ,   A  3;   A  3�   �  3�   �  3;   A  3;      B  , ,   A  4�   A  5M   �  5M   �  4�   A  4�      B  , ,   A  6   A  6�   �  6�   �  6   A  6      B  , ,   A  7s   A  8   �  8   �  7s   A  7s      B  , ,    ;    �  �  �  �  ;    ;      B  , ,    �    M  �  M  �  �    �      B  , ,    	    	�  �  	�  �  	    	      B  , ,    
s      �    �  
s    
s      B  , ,    �    �  �  �  �  �    �      B  , ,    C    �  �  �  �  C    C      B  , ,    �    U  �  U  �  �    �      B  , ,        �  �  �  �            B  , ,    {    %  �  %  �  {    {      B  , ,    �    �  �  �  �  �    �      B  , ,    K    �  �  �  �  K    K      B  , ,    �    ]  �  ]  �  �    �      B  , ,        �  �  �  �            B  , ,    �    -  �  -  �  �    �      B  , ,    �    �  �  �  �  �    �      B  , ,    S    �  �  �  �  S    S      B  , ,    �    e  �  e  �  �    �      B  , ,  �    �  �  S  �  S    �        B  , ,  �  k  �    S    S  k  �  k      B  , ,  �  �  �  }  S  }  S  �  �  �      B  , ,  �  ;  �  �  S  �  S  ;  �  ;      B  , ,  �  �  �  M  S  M  S  �  �  �      B  , ,  �  	  �  	�  S  	�  S  	  �  	      B  , ,  �  
s  �    S    S  
s  �  
s      B  , ,  �  �  �  �  S  �  S  �  �  �      B  , ,  �  C  �  �  S  �  S  C  �  C      B  , ,  �  �  �  U  S  U  S  �  �  �      B  , ,  �    �  �  S  �  S    �        B  , ,  �  {  �  %  S  %  S  {  �  {      B  , ,  �  �  �  �  S  �  S  �  �  �      B  , ,  �  K  �  �  S  �  S  K  �  K      B  , ,  �  �  �  ]  S  ]  S  �  �  �      B  , ,  �    �  �  S  �  S    �        B  , ,  �  �  �  -  S  -  S  �  �  �      B  , ,  �  �  �  �  S  �  S  �  �  �      B  , ,  �  S  �  �  S  �  S  S  �  S      B  , ,  �  �  �  e  S  e  S  �  �  �      B  , ,  
�  
s  
�    O    O  
s  
�  
s      B  , ,  
�  �  
�  �  O  �  O  �  
�  �      B  , ,  
�  C  
�  �  O  �  O  C  
�  C      B  , ,  
�  �  
�  U  O  U  O  �  
�  �      B  , ,   A   �   A  E   �  E   �   �   A   �      B  , ,   A     A  �   �  �   �     A        B  , ,   A  k   A     �     �  k   A  k      B  , ,   A  �   A  }   �  }   �  �   A  �      B  , ,   A  ;   A  �   �  �   �  ;   A  ;      B  , ,   A  �   A  M   �  M   �  �   A  �      B  , ,   A  	   A  	�   �  	�   �  	   A  	      B  , ,   A  
s   A     �     �  
s   A  
s      B  , ,   A  �   A  �   �  �   �  �   A  �      B  , ,   A  C   A  �   �  �   �  C   A  C      B  , ,   A  �   A  U   �  U   �  �   A  �      B  , ,   A     A  �   �  �   �     A        B  , ,   A  {   A  %   �  %   �  {   A  {      B  , ,   A  �   A  �   �  �   �  �   A  �      B  , ,   A  K   A  �   �  �   �  K   A  K      B  , ,   A  �   A  ]   �  ]   �  �   A  �      B  , ,   A     A  �   �  �   �     A        B  , ,   A  �   A  -   �  -   �  �   A  �      B  , ,   A  �   A  �   �  �   �  �   A  �      B  , ,   A  S   A  �   �  �   �  S   A  S      B  , ,   A  �   A  e   �  e   �  �   A  �      B  , ,  
�    
�  �  O  �  O    
�        B  , ,  
�  {  
�  %  O  %  O  {  
�  {      B  , ,  
�  �  
�  �  O  �  O  �  
�  �      B  , ,  
�  K  
�  �  O  �  O  K  
�  K      B  , ,  
�  �  
�  ]  O  ]  O  �  
�  �      B  , ,  
�    
�  �  O  �  O    
�        B  , ,  
�  �  
�  -  O  -  O  �  
�  �      B  , ,  
�  �  
�  �  O  �  O  �  
�  �      B  , ,  
�  S  
�  �  O  �  O  S  
�  S      B  , ,  
�  �  
�  e  O  e  O  �  
�  �      B  , ,  
�  �  
�  }  O  }  O  �  
�  �      B  , ,  
�  ;  
�  �  O  �  O  ;  
�  ;      B  , ,  
�  �  
�  M  O  M  O  �  
�  �      B  , ,  
�  	  
�  	�  O  	�  O  	  
�  	      B  , ,  �   �  �  E  S  E  S   �  �   �      B  , ,     �    E  �  E  �   �     �      B  , ,        �  �  �  �            B  , ,    k      �    �  k    k      B  , ,    �    }  �  }  �  �    �      B  , ,  
�   �  
�  E  O  E  O   �  
�   �      B  , ,  
�    
�  �  O  �  O    
�        B  , ,  
�  k  
�    O    O  k  
�  k      A   ,              u0  �  u0  �                  ]  , ,������������  u�  u  u�  u������������     � 
   % 0� 
   % 0 nfet    B   ,  ,���8  ,  �  �  �  ����8  ,���8      B   ,  	  �  	  �    �    �  	  �      A  , ,            �  �  �  �                 D   ,   #   �   #  9  	  9  	   �   #   �      D   ,     �    9  �  9  �   �     �      D   ,   �  �   �  �  G  �  G  �   �  �      _   ,   �  �   �    !    !  �   �  �      C   ,   A   �   A  M   �  M   �   �   A   �      C   ,  5   �  5  M  �  M  �   �  5   �      C   ,   �      �  �  5  �  5      �         C   ,  �   �  �  M  V  M  V   �  �   �      ^   ,   ����     e  ^  e  ^����   ����      C  , ,   A   �   A  �   �  �   �   �   A   �      C  , ,   A  S   A  �   �  �   �  S   A  S      C  , ,  5   �  5  �  �  �  �   �  5   �      C  , ,  5  S  5  �  �  �  �  S  5  S      C  , ,  ;     ;  �  �  �  �     ;         B  , ,   A   �   A  �   �  �   �   �   A   �      B  , ,   A  S   A  �   �  �   �  S   A  S      B  , ,  5   �  5  �  �  �  �   �  5   �      B  , ,  5  S  5  �  �  �  �  S  5  S      B  , ,  ;     ;  �  �  �  �     ;         B  , ,  �   �  �  �  V  �  V   �  �   �      B  , ,  �  S  �  �  V  �  V  S  �  S      A   ,              �     �                     ]  , ,������������  e    e  ������������     � 
   % 0� 
   % 0 inv_strvd  
  nfet$10     BZ         '�  �   
  
pfet$6    BZ         O  �   
  nfet �  C�      ���c  I      D   ,����  �����  �����  �����  �����  �      D   ,����������   2����   2���������������      D   ,���  p���  h  N�  h  N�  p���  p      D   ,�������c����  ���a  ���a���c�������c      D   ,����  ����  $�����  $�����  ����        D   ,���  p���  h  N�  h  N�  p���  p      D   ,����  ����  $�����  $�����  ����        D   ,���  @���  Z����  Z����  @���  @      D   ,���  )���  -�  N�  -�  N�  )���  )      D   ,  N�  *  N�  -�  N�  -�  N�  *  N�  *      D   ,����  *����  -����  -����  *����  *      C  , ,   �  *   �  *�  @  *�  @  *   �  *      C  , ,   �  +i   �  ,  @  ,  @  +i   �  +i      C  , ,   �  ,�   �  -{  @  -{  @  ,�   �  ,�      C  , ,  '�  *  '�  *�  (�  *�  (�  *  '�  *      C  , ,  )^  *  )^  *�  *  *�  *  *  )^  *      C  , ,  *�  *  *�  *�  +p  *�  +p  *  *�  *      C  , ,  ,.  *  ,.  *�  ,�  *�  ,�  *  ,.  *      C  , ,  -�  *  -�  *�  .@  *�  .@  *  -�  *      C  , ,  .�  *  .�  *�  /�  *�  /�  *  .�  *      C  , ,  0f  *  0f  *�  1  *�  1  *  0f  *      C  , ,  1�  *  1�  *�  2x  *�  2x  *  1�  *      C  , ,  36  *  36  *�  3�  *�  3�  *  36  *      C  , ,  4�  *  4�  *�  5H  *�  5H  *  4�  *      C  , ,  6  *  6  *�  6�  *�  6�  *  6  *      C  , ,  7n  *  7n  *�  8  *�  8  *  7n  *      C  , ,  8�  *  8�  *�  9�  *�  9�  *  8�  *      C  , ,  :>  *  :>  *�  :�  *�  :�  *  :>  *      C  , ,  ;�  *  ;�  *�  <P  *�  <P  *  ;�  *      C  , ,  =  *  =  *�  =�  *�  =�  *  =  *      C  , ,  >v  *  >v  *�  ?   *�  ?   *  >v  *      C  , ,  ?�  *  ?�  *�  @�  *�  @�  *  ?�  *      C  , ,  AF  *  AF  *�  A�  *�  A�  *  AF  *      C  , ,  B�  *  B�  *�  CX  *�  CX  *  B�  *      C  , ,  D  *  D  *�  D�  *�  D�  *  D  *      C  , ,  E~  *  E~  *�  F(  *�  F(  *  E~  *      C  , ,  F�  *  F�  *�  G�  *�  G�  *  F�  *      C  , ,  HN  *  HN  *�  H�  *�  H�  *  HN  *      C  , ,  I�  *  I�  *�  J`  *�  J`  *  I�  *      C  , ,  K  *  K  *�  K�  *�  K�  *  K  *      C  , ,  L�  *  L�  *�  M0  *�  M0  *  L�  *      C  , ,  M�  *  M�  *�  N�  *�  N�  *  M�  *      C  , ,  '�  +i  '�  ,  (�  ,  (�  +i  '�  +i      C  , ,  )^  +i  )^  ,  *  ,  *  +i  )^  +i      C  , ,  *�  +i  *�  ,  +p  ,  +p  +i  *�  +i      C  , ,  ,.  +i  ,.  ,  ,�  ,  ,�  +i  ,.  +i      C  , ,  -�  +i  -�  ,  .@  ,  .@  +i  -�  +i      C  , ,  .�  +i  .�  ,  /�  ,  /�  +i  .�  +i      C  , ,  0f  +i  0f  ,  1  ,  1  +i  0f  +i      C  , ,  1�  +i  1�  ,  2x  ,  2x  +i  1�  +i      C  , ,  36  +i  36  ,  3�  ,  3�  +i  36  +i      C  , ,  4�  +i  4�  ,  5H  ,  5H  +i  4�  +i      C  , ,  6  +i  6  ,  6�  ,  6�  +i  6  +i      C  , ,  7n  +i  7n  ,  8  ,  8  +i  7n  +i      C  , ,  8�  +i  8�  ,  9�  ,  9�  +i  8�  +i      C  , ,  :>  +i  :>  ,  :�  ,  :�  +i  :>  +i      C  , ,  ;�  +i  ;�  ,  <P  ,  <P  +i  ;�  +i      C  , ,  =  +i  =  ,  =�  ,  =�  +i  =  +i      C  , ,  >v  +i  >v  ,  ?   ,  ?   +i  >v  +i      C  , ,  ?�  +i  ?�  ,  @�  ,  @�  +i  ?�  +i      C  , ,  AF  +i  AF  ,  A�  ,  A�  +i  AF  +i      C  , ,  B�  +i  B�  ,  CX  ,  CX  +i  B�  +i      C  , ,  D  +i  D  ,  D�  ,  D�  +i  D  +i      C  , ,  E~  +i  E~  ,  F(  ,  F(  +i  E~  +i      C  , ,  F�  +i  F�  ,  G�  ,  G�  +i  F�  +i      C  , ,  HN  +i  HN  ,  H�  ,  H�  +i  HN  +i      C  , ,  I�  +i  I�  ,  J`  ,  J`  +i  I�  +i      C  , ,  K  +i  K  ,  K�  ,  K�  +i  K  +i      C  , ,  L�  +i  L�  ,  M0  ,  M0  +i  L�  +i      C  , ,  M�  +i  M�  ,  N�  ,  N�  +i  M�  +i      C  , ,  '�  ,�  '�  -{  (�  -{  (�  ,�  '�  ,�      C  , ,  )^  ,�  )^  -{  *  -{  *  ,�  )^  ,�      C  , ,  *�  ,�  *�  -{  +p  -{  +p  ,�  *�  ,�      C  , ,  ,.  ,�  ,.  -{  ,�  -{  ,�  ,�  ,.  ,�      C  , ,  -�  ,�  -�  -{  .@  -{  .@  ,�  -�  ,�      C  , ,  .�  ,�  .�  -{  /�  -{  /�  ,�  .�  ,�      C  , ,  0f  ,�  0f  -{  1  -{  1  ,�  0f  ,�      C  , ,  1�  ,�  1�  -{  2x  -{  2x  ,�  1�  ,�      C  , ,  36  ,�  36  -{  3�  -{  3�  ,�  36  ,�      C  , ,  4�  ,�  4�  -{  5H  -{  5H  ,�  4�  ,�      C  , ,  6  ,�  6  -{  6�  -{  6�  ,�  6  ,�      C  , ,  7n  ,�  7n  -{  8  -{  8  ,�  7n  ,�      C  , ,  8�  ,�  8�  -{  9�  -{  9�  ,�  8�  ,�      C  , ,  :>  ,�  :>  -{  :�  -{  :�  ,�  :>  ,�      C  , ,  ;�  ,�  ;�  -{  <P  -{  <P  ,�  ;�  ,�      C  , ,  =  ,�  =  -{  =�  -{  =�  ,�  =  ,�      C  , ,  >v  ,�  >v  -{  ?   -{  ?   ,�  >v  ,�      C  , ,  ?�  ,�  ?�  -{  @�  -{  @�  ,�  ?�  ,�      C  , ,  AF  ,�  AF  -{  A�  -{  A�  ,�  AF  ,�      C  , ,  B�  ,�  B�  -{  CX  -{  CX  ,�  B�  ,�      C  , ,  D  ,�  D  -{  D�  -{  D�  ,�  D  ,�      C  , ,  E~  ,�  E~  -{  F(  -{  F(  ,�  E~  ,�      C  , ,  F�  ,�  F�  -{  G�  -{  G�  ,�  F�  ,�      C  , ,  HN  ,�  HN  -{  H�  -{  H�  ,�  HN  ,�      C  , ,  I�  ,�  I�  -{  J`  -{  J`  ,�  I�  ,�      C  , ,  K  ,�  K  -{  K�  -{  K�  ,�  K  ,�      C  , ,  L�  ,�  L�  -{  M0  -{  M0  ,�  L�  ,�      C  , ,  M�  ,�  M�  -{  N�  -{  N�  ,�  M�  ,�      C  , ,  >  *  >  *�  �  *�  �  *  >  *      C  , ,  �  *  �  *�  P  *�  P  *  �  *      C  , ,    *    *�  �  *�  �  *    *      C  , ,  v  *  v  *�     *�     *  v  *      C  , ,  �  *  �  *�  �  *�  �  *  �  *      C  , ,  F  *  F  *�  �  *�  �  *  F  *      C  , ,  �  *  �  *�  X  *�  X  *  �  *      C  , ,    *    *�  �  *�  �  *    *      C  , ,  ~  *  ~  *�  (  *�  (  *  ~  *      C  , ,  �  *  �  *�  �  *�  �  *  �  *      C  , ,  N  *  N  *�  �  *�  �  *  N  *      C  , ,  �  *  �  *�  `  *�  `  *  �  *      C  , ,    *    *�  �  *�  �  *    *      C  , ,  �  *  �  *�   0  *�   0  *  �  *      C  , ,   �  *   �  *�  !�  *�  !�  *   �  *      C  , ,  "V  *  "V  *�  #   *�  #   *  "V  *      C  , ,  #�  *  #�  *�  $h  *�  $h  *  #�  *      C  , ,  %&  *  %&  *�  %�  *�  %�  *  %&  *      C  , ,  &�  *  &�  *�  '8  *�  '8  *  &�  *      C  , ,  �  *  �  *�  x  *�  x  *  �  *      C  , ,  6  *  6  *�  �  *�  �  *  6  *      C  , ,  �  *  �  *�  H  *�  H  *  �  *      C  , ,  �  *  �  *�  �  *�  �  *  �  *      C  , ,  �  +i  �  ,  �  ,  �  +i  �  +i      C  , ,  f  +i  f  ,    ,    +i  f  +i      C  , ,  f  *  f  *�    *�    *  f  *      C  , ,  �  ,�  �  -{  �  -{  �  ,�  �  ,�      C  , ,  f  ,�  f  -{    -{    ,�  f  ,�      C  , ,  �  ,�  �  -{  x  -{  x  ,�  �  ,�      C  , ,  6  ,�  6  -{  �  -{  �  ,�  6  ,�      C  , ,  �  ,�  �  -{  H  -{  H  ,�  �  ,�      C  , ,  	  ,�  	  -{  	�  -{  	�  ,�  	  ,�      C  , ,  
n  ,�  
n  -{    -{    ,�  
n  ,�      C  , ,  �  ,�  �  -{  �  -{  �  ,�  �  ,�      C  , ,  >  ,�  >  -{  �  -{  �  ,�  >  ,�      C  , ,  �  ,�  �  -{  P  -{  P  ,�  �  ,�      C  , ,    ,�    -{  �  -{  �  ,�    ,�      C  , ,  v  ,�  v  -{     -{     ,�  v  ,�      C  , ,  �  ,�  �  -{  �  -{  �  ,�  �  ,�      C  , ,  F  ,�  F  -{  �  -{  �  ,�  F  ,�      C  , ,  �  ,�  �  -{  X  -{  X  ,�  �  ,�      C  , ,    ,�    -{  �  -{  �  ,�    ,�      C  , ,  ~  ,�  ~  -{  (  -{  (  ,�  ~  ,�      C  , ,  �  ,�  �  -{  �  -{  �  ,�  �  ,�      C  , ,  N  ,�  N  -{  �  -{  �  ,�  N  ,�      C  , ,  �  ,�  �  -{  `  -{  `  ,�  �  ,�      C  , ,    ,�    -{  �  -{  �  ,�    ,�      C  , ,  �  ,�  �  -{   0  -{   0  ,�  �  ,�      C  , ,   �  ,�   �  -{  !�  -{  !�  ,�   �  ,�      C  , ,  "V  ,�  "V  -{  #   -{  #   ,�  "V  ,�      C  , ,  #�  ,�  #�  -{  $h  -{  $h  ,�  #�  ,�      C  , ,  %&  ,�  %&  -{  %�  -{  %�  ,�  %&  ,�      C  , ,  &�  ,�  &�  -{  '8  -{  '8  ,�  &�  ,�      C  , ,  �  +i  �  ,  x  ,  x  +i  �  +i      C  , ,  6  +i  6  ,  �  ,  �  +i  6  +i      C  , ,  �  +i  �  ,  H  ,  H  +i  �  +i      C  , ,  	  +i  	  ,  	�  ,  	�  +i  	  +i      C  , ,  
n  +i  
n  ,    ,    +i  
n  +i      C  , ,  �  +i  �  ,  �  ,  �  +i  �  +i      C  , ,  >  +i  >  ,  �  ,  �  +i  >  +i      C  , ,  �  +i  �  ,  P  ,  P  +i  �  +i      C  , ,    +i    ,  �  ,  �  +i    +i      C  , ,  v  +i  v  ,     ,     +i  v  +i      C  , ,  �  +i  �  ,  �  ,  �  +i  �  +i      C  , ,  F  +i  F  ,  �  ,  �  +i  F  +i      C  , ,  �  +i  �  ,  X  ,  X  +i  �  +i      C  , ,    +i    ,  �  ,  �  +i    +i      C  , ,  ~  +i  ~  ,  (  ,  (  +i  ~  +i      C  , ,  �  +i  �  ,  �  ,  �  +i  �  +i      C  , ,  N  +i  N  ,  �  ,  �  +i  N  +i      C  , ,  �  +i  �  ,  `  ,  `  +i  �  +i      C  , ,    +i    ,  �  ,  �  +i    +i      C  , ,  �  +i  �  ,   0  ,   0  +i  �  +i      C  , ,   �  +i   �  ,  !�  ,  !�  +i   �  +i      C  , ,  "V  +i  "V  ,  #   ,  #   +i  "V  +i      C  , ,  #�  +i  #�  ,  $h  ,  $h  +i  #�  +i      C  , ,  %&  +i  %&  ,  %�  ,  %�  +i  %&  +i      C  , ,  &�  +i  &�  ,  '8  ,  '8  +i  &�  +i      C  , ,  	  *  	  *�  	�  *�  	�  *  	  *      C  , ,  
n  *  
n  *�    *�    *  
n  *      C  , ,  �  *  �  *�  �  *�  �  *  �  *      C  , ,��ڞ  +i��ڞ  ,���H  ,���H  +i��ڞ  +i      C  , ,���  +i���  ,��ܰ  ,��ܰ  +i���  +i      C  , ,���n  +i���n  ,���  ,���  +i���n  +i      C  , ,����  +i����  ,��߀  ,��߀  +i����  +i      C  , ,���>  +i���>  ,����  ,����  +i���>  +i      C  , ,���  +i���  ,���P  ,���P  +i���  +i      C  , ,���  +i���  ,���  ,���  +i���  +i      C  , ,���v  +i���v  ,���   ,���   +i���v  +i      C  , ,����  +i����  ,���  ,���  +i����  +i      C  , ,���F  +i���F  ,����  ,����  +i���F  +i      C  , ,���  +i���  ,���X  ,���X  +i���  +i      C  , ,���  +i���  ,����  ,����  +i���  +i      C  , ,���~  +i���~  ,���(  ,���(  +i���~  +i      C  , ,����  +i����  ,���  ,���  +i����  +i      C  , ,���N  +i���N  ,����  ,����  +i���N  +i      C  , ,���  +i���  ,���`  ,���`  +i���  +i      C  , ,���  +i���  ,����  ,����  +i���  +i      C  , ,���  +i���  ,���0  ,���0  +i���  +i      C  , ,����  +i����  ,����  ,����  +i����  +i      C  , ,���V  +i���V  ,���   ,���   +i���V  +i      C  , ,����  +i����  ,���h  ,���h  +i����  +i      C  , ,���&  +i���&  ,����  ,����  +i���&  +i      C  , ,����  +i����  ,���8  ,���8  +i����  +i      C  , ,����  +i����  ,����  ,����  +i����  +i      C  , ,���^  +i���^  ,���  ,���  +i���^  +i      C  , ,����  +i����  ,���p  ,���p  +i����  +i      C  , ,���.  +i���.  ,����  ,����  +i���.  +i      C  , ,��ڞ  *��ڞ  *����H  *����H  *��ڞ  *      C  , ,���  *���  *���ܰ  *���ܰ  *���  *      C  , ,���n  *���n  *����  *����  *���n  *      C  , ,����  *����  *���߀  *���߀  *����  *      C  , ,���>  *���>  *�����  *�����  *���>  *      C  , ,���  *���  *����P  *����P  *���  *      C  , ,���  *���  *����  *����  *���  *      C  , ,���v  *���v  *����   *����   *���v  *      C  , ,����  *����  *����  *����  *����  *      C  , ,���F  *���F  *�����  *�����  *���F  *      C  , ,���  *���  *����X  *����X  *���  *      C  , ,���  *���  *�����  *�����  *���  *      C  , ,���~  *���~  *����(  *����(  *���~  *      C  , ,����  *����  *����  *����  *����  *      C  , ,���N  *���N  *�����  *�����  *���N  *      C  , ,���  *���  *����`  *����`  *���  *      C  , ,���  *���  *�����  *�����  *���  *      C  , ,���  *���  *����0  *����0  *���  *      C  , ,����  *����  *�����  *�����  *����  *      C  , ,���V  *���V  *����   *����   *���V  *      C  , ,����  *����  *����h  *����h  *����  *      C  , ,���&  *���&  *�����  *�����  *���&  *      C  , ,����  *����  *����8  *����8  *����  *      C  , ,����  *����  *�����  *�����  *����  *      C  , ,���^  *���^  *����  *����  *���^  *      C  , ,����  *����  *����p  *����p  *����  *      C  , ,���.  *���.  *�����  *�����  *���.  *      C  , ,��ڞ  ,���ڞ  -{���H  -{���H  ,���ڞ  ,�      C  , ,���  ,����  -{��ܰ  -{��ܰ  ,����  ,�      C  , ,���n  ,����n  -{���  -{���  ,����n  ,�      C  , ,����  ,�����  -{��߀  -{��߀  ,�����  ,�      C  , ,���>  ,����>  -{����  -{����  ,����>  ,�      C  , ,���  ,����  -{���P  -{���P  ,����  ,�      C  , ,���  ,����  -{���  -{���  ,����  ,�      C  , ,���v  ,����v  -{���   -{���   ,����v  ,�      C  , ,����  ,�����  -{���  -{���  ,�����  ,�      C  , ,���F  ,����F  -{����  -{����  ,����F  ,�      C  , ,���  ,����  -{���X  -{���X  ,����  ,�      C  , ,���  ,����  -{����  -{����  ,����  ,�      C  , ,���~  ,����~  -{���(  -{���(  ,����~  ,�      C  , ,����  ,�����  -{���  -{���  ,�����  ,�      C  , ,���N  ,����N  -{����  -{����  ,����N  ,�      C  , ,���  ,����  -{���`  -{���`  ,����  ,�      C  , ,���  ,����  -{����  -{����  ,����  ,�      C  , ,���  ,����  -{���0  -{���0  ,����  ,�      C  , ,����  ,�����  -{����  -{����  ,�����  ,�      C  , ,���V  ,����V  -{���   -{���   ,����V  ,�      C  , ,����  ,�����  -{���h  -{���h  ,�����  ,�      C  , ,���&  ,����&  -{����  -{����  ,����&  ,�      C  , ,����  ,�����  -{���8  -{���8  ,�����  ,�      C  , ,����  ,�����  -{����  -{����  ,�����  ,�      C  , ,���^  ,����^  -{���  -{���  ,����^  ,�      C  , ,����  ,�����  -{���p  -{���p  ,�����  ,�      C  , ,���.  ,����.  -{����  -{����  ,����.  ,�      C  , ,���F  +i���F  ,����  ,����  +i���F  +i      C  , ,����  +i����  ,���X  ,���X  +i����  +i      C  , ,���  +i���  ,����  ,����  +i���  +i      C  , ,���~  +i���~  ,���(  ,���(  +i���~  +i      C  , ,����  +i����  ,����  ,����  +i����  +i      C  , ,���N  +i���N  ,����  ,����  +i���N  +i      C  , ,��¶  +i��¶  ,���`  ,���`  +i��¶  +i      C  , ,���  +i���  ,����  ,����  +i���  +i      C  , ,��ņ  +i��ņ  ,���0  ,���0  +i��ņ  +i      C  , ,����  +i����  ,��ǘ  ,��ǘ  +i����  +i      C  , ,���V  +i���V  ,���   ,���   +i���V  +i      C  , ,��ɾ  +i��ɾ  ,���h  ,���h  +i��ɾ  +i      C  , ,���&  +i���&  ,����  ,����  +i���&  +i      C  , ,��̎  +i��̎  ,���8  ,���8  +i��̎  +i      C  , ,����  +i����  ,��Π  ,��Π  +i����  +i      C  , ,���^  +i���^  ,���  ,���  +i���^  +i      C  , ,����  +i����  ,���p  ,���p  +i����  +i      C  , ,���.  +i���.  ,����  ,����  +i���.  +i      C  , ,��Ӗ  +i��Ӗ  ,���@  ,���@  +i��Ӗ  +i      C  , ,����  +i����  ,��ը  ,��ը  +i����  +i      C  , ,���f  +i���f  ,���  ,���  +i���f  +i      C  , ,����  +i����  ,���x  ,���x  +i����  +i      C  , ,���6  +i���6  ,����  ,����  +i���6  +i      C  , ,���  +i���  ,����  ,����  +i���  +i      C  , ,���  *���  *�����  *�����  *���  *      C  , ,���>  *���>  *�����  *�����  *���>  *      C  , ,����  *����  *����P  *����P  *����  *      C  , ,����  +i����  ,���P  ,���P  +i����  +i      C  , ,����  ,�����  -{���P  -{���P  ,�����  ,�      C  , ,���  ,����  -{����  -{����  ,����  ,�      C  , ,���v  ,����v  -{���   -{���   ,����v  ,�      C  , ,����  ,�����  -{����  -{����  ,�����  ,�      C  , ,���F  ,����F  -{����  -{����  ,����F  ,�      C  , ,����  ,�����  -{���X  -{���X  ,�����  ,�      C  , ,���  ,����  -{����  -{����  ,����  ,�      C  , ,���~  ,����~  -{���(  -{���(  ,����~  ,�      C  , ,����  ,�����  -{����  -{����  ,�����  ,�      C  , ,���N  ,����N  -{����  -{����  ,����N  ,�      C  , ,��¶  ,���¶  -{���`  -{���`  ,���¶  ,�      C  , ,���  ,����  -{����  -{����  ,����  ,�      C  , ,��ņ  ,���ņ  -{���0  -{���0  ,���ņ  ,�      C  , ,����  ,�����  -{��ǘ  -{��ǘ  ,�����  ,�      C  , ,���V  ,����V  -{���   -{���   ,����V  ,�      C  , ,��ɾ  ,���ɾ  -{���h  -{���h  ,���ɾ  ,�      C  , ,���&  ,����&  -{����  -{����  ,����&  ,�      C  , ,��̎  ,���̎  -{���8  -{���8  ,���̎  ,�      C  , ,����  ,�����  -{��Π  -{��Π  ,�����  ,�      C  , ,���^  ,����^  -{���  -{���  ,����^  ,�      C  , ,����  ,�����  -{���p  -{���p  ,�����  ,�      C  , ,���.  ,����.  -{����  -{����  ,����.  ,�      C  , ,��Ӗ  ,���Ӗ  -{���@  -{���@  ,���Ӗ  ,�      C  , ,����  ,�����  -{��ը  -{��ը  ,�����  ,�      C  , ,���f  ,����f  -{���  -{���  ,����f  ,�      C  , ,����  ,�����  -{���x  -{���x  ,�����  ,�      C  , ,���6  ,����6  -{����  -{����  ,����6  ,�      C  , ,���v  *���v  *����   *����   *���v  *      C  , ,����  *����  *�����  *�����  *����  *      C  , ,���F  *���F  *�����  *�����  *���F  *      C  , ,����  *����  *����X  *����X  *����  *      C  , ,���  *���  *�����  *�����  *���  *      C  , ,���~  *���~  *����(  *����(  *���~  *      C  , ,����  *����  *�����  *�����  *����  *      C  , ,���N  *���N  *�����  *�����  *���N  *      C  , ,��¶  *��¶  *����`  *����`  *��¶  *      C  , ,���  *���  *�����  *�����  *���  *      C  , ,��ņ  *��ņ  *����0  *����0  *��ņ  *      C  , ,����  *����  *���ǘ  *���ǘ  *����  *      C  , ,���V  *���V  *����   *����   *���V  *      C  , ,��ɾ  *��ɾ  *����h  *����h  *��ɾ  *      C  , ,���&  *���&  *�����  *�����  *���&  *      C  , ,��̎  *��̎  *����8  *����8  *��̎  *      C  , ,����  *����  *���Π  *���Π  *����  *      C  , ,���^  *���^  *����  *����  *���^  *      C  , ,����  *����  *����p  *����p  *����  *      C  , ,���.  *���.  *�����  *�����  *���.  *      C  , ,��Ӗ  *��Ӗ  *����@  *����@  *��Ӗ  *      C  , ,����  *����  *���ը  *���ը  *����  *      C  , ,���f  *���f  *����  *����  *���f  *      C  , ,����  *����  *����x  *����x  *����  *      C  , ,���6  *���6  *�����  *�����  *���6  *      C  , ,���v  +i���v  ,���   ,���   +i���v  +i      C  , ,����  +i����  ,����  ,����  +i����  +i      C  , ,���>  +i���>  ,����  ,����  +i���>  +i      C  , ,���>  ,����>  -{����  -{����  ,����>  ,�      C  , ,�������������������x�������x������������      C  , ,���f�������f���������������������f����      D   ,���  p���  h  N�  h  N�  p���  p      D   ,����  ����  $�����  $�����  ����        D   ,������������  ����4  ����4������������      D     ���   � CTRL      D       N  { OUT       D     ����  � OUT       D       z  � OUT       D       +�  � OUT       D     ��װ  k OUT       D     ����  $T IN      D     ����  � IN      D     ����  � IN      D     ����  � IN      D     ����  J IN      D  , ,   �  *   �  *�  6  *�  6  *   �  *      D  , ,   �  +s   �  ,	  6  ,	  6  +s   �  +s      D  , ,   �  ,�   �  -q  6  -q  6  ,�   �  ,�      D  , ,  0p  +s  0p  ,	  1  ,	  1  +s  0p  +s      D  , ,  1�  +s  1�  ,	  2n  ,	  2n  +s  1�  +s      D  , ,  3@  +s  3@  ,	  3�  ,	  3�  +s  3@  +s      D  , ,  B�  ,�  B�  -q  CN  -q  CN  ,�  B�  ,�      D  , ,  4�  +s  4�  ,	  5>  ,	  5>  +s  4�  +s      D  , ,  D   ,�  D   -q  D�  -q  D�  ,�  D   ,�      D  , ,  6  +s  6  ,	  6�  ,	  6�  +s  6  +s      D  , ,  E�  ,�  E�  -q  F  -q  F  ,�  E�  ,�      D  , ,  7x  +s  7x  ,	  8  ,	  8  +s  7x  +s      D  , ,  F�  ,�  F�  -q  G�  -q  G�  ,�  F�  ,�      D  , ,  8�  +s  8�  ,	  9v  ,	  9v  +s  8�  +s      D  , ,  HX  ,�  HX  -q  H�  -q  H�  ,�  HX  ,�      D  , ,  :H  +s  :H  ,	  :�  ,	  :�  +s  :H  +s      D  , ,  I�  ,�  I�  -q  JV  -q  JV  ,�  I�  ,�      D  , ,  ;�  +s  ;�  ,	  <F  ,	  <F  +s  ;�  +s      D  , ,  K(  ,�  K(  -q  K�  -q  K�  ,�  K(  ,�      D  , ,  =  +s  =  ,	  =�  ,	  =�  +s  =  +s      D  , ,  L�  ,�  L�  -q  M&  -q  M&  ,�  L�  ,�      D  , ,  >�  +s  >�  ,	  ?  ,	  ?  +s  >�  +s      D  , ,  M�  ,�  M�  -q  N�  -q  N�  ,�  M�  ,�      D  , ,  ?�  +s  ?�  ,	  @~  ,	  @~  +s  ?�  +s      D  , ,  (   *  (   *�  (�  *�  (�  *  (   *      D  , ,  AP  +s  AP  ,	  A�  ,	  A�  +s  AP  +s      D  , ,  )h  *  )h  *�  )�  *�  )�  *  )h  *      D  , ,  B�  +s  B�  ,	  CN  ,	  CN  +s  B�  +s      D  , ,  *�  *  *�  *�  +f  *�  +f  *  *�  *      D  , ,  D   +s  D   ,	  D�  ,	  D�  +s  D   +s      D  , ,  ,8  *  ,8  *�  ,�  *�  ,�  *  ,8  *      D  , ,  E�  +s  E�  ,	  F  ,	  F  +s  E�  +s      D  , ,  -�  *  -�  *�  .6  *�  .6  *  -�  *      D  , ,  F�  +s  F�  ,	  G�  ,	  G�  +s  F�  +s      D  , ,  /  *  /  *�  /�  *�  /�  *  /  *      D  , ,  HX  +s  HX  ,	  H�  ,	  H�  +s  HX  +s      D  , ,  0p  *  0p  *�  1  *�  1  *  0p  *      D  , ,  I�  +s  I�  ,	  JV  ,	  JV  +s  I�  +s      D  , ,  1�  *  1�  *�  2n  *�  2n  *  1�  *      D  , ,  K(  +s  K(  ,	  K�  ,	  K�  +s  K(  +s      D  , ,  3@  *  3@  *�  3�  *�  3�  *  3@  *      D  , ,  L�  +s  L�  ,	  M&  ,	  M&  +s  L�  +s      D  , ,  4�  *  4�  *�  5>  *�  5>  *  4�  *      D  , ,  M�  +s  M�  ,	  N�  ,	  N�  +s  M�  +s      D  , ,  6  *  6  *�  6�  *�  6�  *  6  *      D  , ,  (   ,�  (   -q  (�  -q  (�  ,�  (   ,�      D  , ,  7x  *  7x  *�  8  *�  8  *  7x  *      D  , ,  )h  ,�  )h  -q  )�  -q  )�  ,�  )h  ,�      D  , ,  8�  *  8�  *�  9v  *�  9v  *  8�  *      D  , ,  *�  ,�  *�  -q  +f  -q  +f  ,�  *�  ,�      D  , ,  :H  *  :H  *�  :�  *�  :�  *  :H  *      D  , ,  ,8  ,�  ,8  -q  ,�  -q  ,�  ,�  ,8  ,�      D  , ,  ;�  *  ;�  *�  <F  *�  <F  *  ;�  *      D  , ,  -�  ,�  -�  -q  .6  -q  .6  ,�  -�  ,�      D  , ,  =  *  =  *�  =�  *�  =�  *  =  *      D  , ,  /  ,�  /  -q  /�  -q  /�  ,�  /  ,�      D  , ,  >�  *  >�  *�  ?  *�  ?  *  >�  *      D  , ,  0p  ,�  0p  -q  1  -q  1  ,�  0p  ,�      D  , ,  1�  ,�  1�  -q  2n  -q  2n  ,�  1�  ,�      D  , ,  ?�  *  ?�  *�  @~  *�  @~  *  ?�  *      D  , ,  3@  ,�  3@  -q  3�  -q  3�  ,�  3@  ,�      D  , ,  AP  *  AP  *�  A�  *�  A�  *  AP  *      D  , ,  B�  *  B�  *�  CN  *�  CN  *  B�  *      D  , ,  4�  ,�  4�  -q  5>  -q  5>  ,�  4�  ,�      D  , ,  D   *  D   *�  D�  *�  D�  *  D   *      D  , ,  E�  *  E�  *�  F  *�  F  *  E�  *      D  , ,  6  ,�  6  -q  6�  -q  6�  ,�  6  ,�      D  , ,  F�  *  F�  *�  G�  *�  G�  *  F�  *      D  , ,  HX  *  HX  *�  H�  *�  H�  *  HX  *      D  , ,  7x  ,�  7x  -q  8  -q  8  ,�  7x  ,�      D  , ,  I�  *  I�  *�  JV  *�  JV  *  I�  *      D  , ,  K(  *  K(  *�  K�  *�  K�  *  K(  *      D  , ,  8�  ,�  8�  -q  9v  -q  9v  ,�  8�  ,�      D  , ,  L�  *  L�  *�  M&  *�  M&  *  L�  *      D  , ,  M�  *  M�  *�  N�  *�  N�  *  M�  *      D  , ,  :H  ,�  :H  -q  :�  -q  :�  ,�  :H  ,�      D  , ,  ;�  ,�  ;�  -q  <F  -q  <F  ,�  ;�  ,�      D  , ,  =  ,�  =  -q  =�  -q  =�  ,�  =  ,�      D  , ,  >�  ,�  >�  -q  ?  -q  ?  ,�  >�  ,�      D  , ,  ?�  ,�  ?�  -q  @~  -q  @~  ,�  ?�  ,�      D  , ,  AP  ,�  AP  -q  A�  -q  A�  ,�  AP  ,�      D  , ,  (   +s  (   ,	  (�  ,	  (�  +s  (   +s      D  , ,  )h  +s  )h  ,	  )�  ,	  )�  +s  )h  +s      D  , ,  *�  +s  *�  ,	  +f  ,	  +f  +s  *�  +s      D  , ,  ,8  +s  ,8  ,	  ,�  ,	  ,�  +s  ,8  +s      D  , ,  -�  +s  -�  ,	  .6  ,	  .6  +s  -�  +s      D  , ,  /  +s  /  ,	  /�  ,	  /�  +s  /  +s      D  , ,  	  +s  	  ,	  	�  ,	  	�  +s  	  +s      D  , ,  
x  +s  
x  ,	    ,	    +s  
x  +s      D  , ,  �  +s  �  ,	  v  ,	  v  +s  �  +s      D  , ,  H  +s  H  ,	  �  ,	  �  +s  H  +s      D  , ,  �  +s  �  ,	  F  ,	  F  +s  �  +s      D  , ,    +s    ,	  �  ,	  �  +s    +s      D  , ,  �  +s  �  ,	    ,	    +s  �  +s      D  , ,  �  +s  �  ,	  ~  ,	  ~  +s  �  +s      D  , ,  P  +s  P  ,	  �  ,	  �  +s  P  +s      D  , ,  �  +s  �  ,	  n  ,	  n  +s  �  +s      D  , ,  @  +s  @  ,	  �  ,	  �  +s  @  +s      D  , ,  �  +s  �  ,	  >  ,	  >  +s  �  +s      D  , ,  &�  *  &�  *�  '.  *�  '.  *  &�  *      D  , ,  &�  ,�  &�  -q  '.  -q  '.  ,�  &�  ,�      D  , ,  p  ,�  p  -q    -q    ,�  p  ,�      D  , ,  �  ,�  �  -q  v  -q  v  ,�  �  ,�      D  , ,  H  ,�  H  -q  �  -q  �  ,�  H  ,�      D  , ,  �  ,�  �  -q  n  -q  n  ,�  �  ,�      D  , ,  �  ,�  �  -q  F  -q  F  ,�  �  ,�      D  , ,    ,�    -q  �  -q  �  ,�    ,�      D  , ,  @  ,�  @  -q  �  -q  �  ,�  @  ,�      D  , ,  �  ,�  �  -q    -q    ,�  �  ,�      D  , ,  �  ,�  �  -q  ~  -q  ~  ,�  �  ,�      D  , ,  �  ,�  �  -q  >  -q  >  ,�  �  ,�      D  , ,  P  ,�  P  -q  �  -q  �  ,�  P  ,�      D  , ,  �  ,�  �  -q  N  -q  N  ,�  �  ,�      D  , ,  	  ,�  	  -q  	�  -q  	�  ,�  	  ,�      D  , ,     ,�     -q  �  -q  �  ,�     ,�      D  , ,  �  ,�  �  -q    -q    ,�  �  ,�      D  , ,  
x  ,�  
x  -q    -q    ,�  
x  ,�      D  , ,     +s     ,	  �  ,	  �  +s     +s      D  , ,    *    *�  �  *�  �  *    *      D  , ,  p  *  p  *�    *�    *  p  *      D  , ,  �  *  �  *�  n  *�  n  *  �  *      D  , ,  @  *  @  *�  �  *�  �  *  @  *      D  , ,  �  *  �  *�  >  *�  >  *  �  *      D  , ,  	  *  	  *�  	�  *�  	�  *  	  *      D  , ,  
x  *  
x  *�    *�    *  
x  *      D  , ,  �  *  �  *�  v  *�  v  *  �  *      D  , ,  H  *  H  *�  �  *�  �  *  H  *      D  , ,  �  *  �  *�  F  *�  F  *  �  *      D  , ,    *    *�  �  *�  �  *    *      D  , ,  �  *  �  *�    *�    *  �  *      D  , ,  �  *  �  *�  ~  *�  ~  *  �  *      D  , ,  P  *  P  *�  �  *�  �  *  P  *      D  , ,  �  *  �  *�  N  *�  N  *  �  *      D  , ,     *     *�  �  *�  �  *     *      D  , ,  �  *  �  *�    *�    *  �  *      D  , ,  �  *  �  *�  �  *�  �  *  �  *      D  , ,  X  *  X  *�  �  *�  �  *  X  *      D  , ,  �  *  �  *�  V  *�  V  *  �  *      D  , ,  (  *  (  *�  �  *�  �  *  (  *      D  , ,  �  *  �  *�   &  *�   &  *  �  *      D  , ,   �  *   �  *�  !�  *�  !�  *   �  *      D  , ,  "`  *  "`  *�  "�  *�  "�  *  "`  *      D  , ,  #�  *  #�  *�  $^  *�  $^  *  #�  *      D  , ,  %0  *  %0  *�  %�  *�  %�  *  %0  *      D  , ,  �  +s  �  ,	    ,	    +s  �  +s      D  , ,  �  ,�  �  -q  �  -q  �  ,�  �  ,�      D  , ,  X  ,�  X  -q  �  -q  �  ,�  X  ,�      D  , ,  �  ,�  �  -q  V  -q  V  ,�  �  ,�      D  , ,  (  ,�  (  -q  �  -q  �  ,�  (  ,�      D  , ,  �  ,�  �  -q   &  -q   &  ,�  �  ,�      D  , ,   �  ,�   �  -q  !�  -q  !�  ,�   �  ,�      D  , ,  "`  ,�  "`  -q  "�  -q  "�  ,�  "`  ,�      D  , ,  #�  ,�  #�  -q  $^  -q  $^  ,�  #�  ,�      D  , ,  %0  ,�  %0  -q  %�  -q  %�  ,�  %0  ,�      D  , ,    +s    ,	  �  ,	  �  +s    +s      D  , ,  %0  +s  %0  ,	  %�  ,	  %�  +s  %0  +s      D  , ,  p  +s  p  ,	    ,	    +s  p  +s      D  , ,  �  +s  �  ,	  �  ,	  �  +s  �  +s      D  , ,  X  +s  X  ,	  �  ,	  �  +s  X  +s      D  , ,  �  +s  �  ,	  V  ,	  V  +s  �  +s      D  , ,  (  +s  (  ,	  �  ,	  �  +s  (  +s      D  , ,  �  +s  �  ,	   &  ,	   &  +s  �  +s      D  , ,   �  +s   �  ,	  !�  ,	  !�  +s   �  +s      D  , ,  "`  +s  "`  ,	  "�  ,	  "�  +s  "`  +s      D  , ,  #�  +s  #�  ,	  $^  ,	  $^  +s  #�  +s      D  , ,  �  +s  �  ,	  N  ,	  N  +s  �  +s      D  , ,    ,�    -q  �  -q  �  ,�    ,�      D  , ,  &�  +s  &�  ,	  '.  ,	  '.  +s  &�  +s      D  , ,���8  +s���8  ,	����  ,	����  +s���8  +s      D  , ,���8  *���8  *�����  *�����  *���8  *      D  , ,���8  ,����8  -q����  -q����  ,����8  ,�      D  , ,���  ,����  -q���  -q���  ,����  ,�      D  , ,���  ,����  -q���  -q���  ,����  ,�      D  , ,����  ,�����  -q���~  -q���~  ,�����  ,�      D  , ,���P  ,����P  -q����  -q����  ,����P  ,�      D  , ,���  ,����  -q���N  -q���N  ,����  ,�      D  , ,���   ,����   -q���  -q���  ,����   ,�      D  , ,���  ,����  -q���  -q���  ,����  ,�      D  , ,����  ,�����  -q���  -q���  ,�����  ,�      D  , ,���X  ,����X  -q����  -q����  ,����X  ,�      D  , ,����  ,�����  -q���V  -q���V  ,�����  ,�      D  , ,���(  ,����(  -q���  -q���  ,����(  ,�      D  , ,���  ,����  -q���&  -q���&  ,����  ,�      D  , ,����  ,�����  -q���  -q���  ,�����  ,�      D  , ,���`  ,����`  -q����  -q����  ,����`  ,�      D  , ,����  ,�����  -q���^  -q���^  ,�����  ,�      D  , ,���0  ,����0  -q����  -q����  ,����0  ,�      D  , ,����  ,�����  -q���.  -q���.  ,�����  ,�      D  , ,���   ,����   -q����  -q����  ,����   ,�      D  , ,���h  ,����h  -q����  -q����  ,����h  ,�      D  , ,����  ,�����  -q���f  -q���f  ,�����  ,�      D  , ,���  *���  *���ܦ  *���ܦ  *���  *      D  , ,��ڨ  +s��ڨ  ,	���>  ,	���>  +s��ڨ  +s      D  , ,���  +s���  ,	��ܦ  ,	��ܦ  +s���  +s      D  , ,���x  +s���x  ,	���  ,	���  +s���x  +s      D  , ,����  +s����  ,	���v  ,	���v  +s����  +s      D  , ,���H  +s���H  ,	����  ,	����  +s���H  +s      D  , ,���  +s���  ,	���F  ,	���F  +s���  +s      D  , ,���  +s���  ,	���  ,	���  +s���  +s      D  , ,���  +s���  ,	���  ,	���  +s���  +s      D  , ,����  +s����  ,	���~  ,	���~  +s����  +s      D  , ,���P  +s���P  ,	����  ,	����  +s���P  +s      D  , ,���  +s���  ,	���N  ,	���N  +s���  +s      D  , ,���   +s���   ,	���  ,	���  +s���   +s      D  , ,���  +s���  ,	���  ,	���  +s���  +s      D  , ,����  +s����  ,	���  ,	���  +s����  +s      D  , ,���X  +s���X  ,	����  ,	����  +s���X  +s      D  , ,����  +s����  ,	���V  ,	���V  +s����  +s      D  , ,���(  +s���(  ,	���  ,	���  +s���(  +s      D  , ,���  +s���  ,	���&  ,	���&  +s���  +s      D  , ,����  +s����  ,	���  ,	���  +s����  +s      D  , ,���`  +s���`  ,	����  ,	����  +s���`  +s      D  , ,����  +s����  ,	���^  ,	���^  +s����  +s      D  , ,���0  +s���0  ,	����  ,	����  +s���0  +s      D  , ,����  +s����  ,	���.  ,	���.  +s����  +s      D  , ,���   +s���   ,	����  ,	����  +s���   +s      D  , ,���h  +s���h  ,	����  ,	����  +s���h  +s      D  , ,����  +s����  ,	���f  ,	���f  +s����  +s      D  , ,���x  *���x  *����  *����  *���x  *      D  , ,����  *����  *����v  *����v  *����  *      D  , ,���H  *���H  *�����  *�����  *���H  *      D  , ,���  *���  *����F  *����F  *���  *      D  , ,���  *���  *����  *����  *���  *      D  , ,���  *���  *����  *����  *���  *      D  , ,����  *����  *����~  *����~  *����  *      D  , ,���P  *���P  *�����  *�����  *���P  *      D  , ,���  *���  *����N  *����N  *���  *      D  , ,���   *���   *����  *����  *���   *      D  , ,���  *���  *����  *����  *���  *      D  , ,����  *����  *����  *����  *����  *      D  , ,���X  *���X  *�����  *�����  *���X  *      D  , ,����  *����  *����V  *����V  *����  *      D  , ,���(  *���(  *����  *����  *���(  *      D  , ,���  *���  *����&  *����&  *���  *      D  , ,����  *����  *����  *����  *����  *      D  , ,���`  *���`  *�����  *�����  *���`  *      D  , ,����  *����  *����^  *����^  *����  *      D  , ,���0  *���0  *�����  *�����  *���0  *      D  , ,��ڨ  ,���ڨ  -q���>  -q���>  ,���ڨ  ,�      D  , ,����  *����  *����.  *����.  *����  *      D  , ,���  ,����  -q��ܦ  -q��ܦ  ,����  ,�      D  , ,���   *���   *�����  *�����  *���   *      D  , ,���x  ,����x  -q���  -q���  ,����x  ,�      D  , ,���h  *���h  *�����  *�����  *���h  *      D  , ,����  ,�����  -q���v  -q���v  ,�����  ,�      D  , ,����  *����  *����f  *����f  *����  *      D  , ,���H  ,����H  -q����  -q����  ,����H  ,�      D  , ,��ڨ  *��ڨ  *����>  *����>  *��ڨ  *      D  , ,���  ,����  -q���F  -q���F  ,����  ,�      D  , ,����  *����  *����n  *����n  *����  *      D  , ,����  +s����  ,	���n  ,	���n  +s����  +s      D  , ,���@  *���@  *�����  *�����  *���@  *      D  , ,���@  ,����@  -q����  -q����  ,����@  ,�      D  , ,���@  +s���@  ,	����  ,	����  +s���@  +s      D  , ,����  ,�����  -q���n  -q���n  ,�����  ,�      D  , ,����  ,�����  -q���  -q���  ,�����  ,�      D  , ,���  *���  *�����  *�����  *���  *      D  , ,���   +s���   ,	����  ,	����  +s���   +s      D  , ,���0  ,����0  -q����  -q����  ,����0  ,�      D  , ,����  +s����  ,	���  ,	���  +s����  +s      D  , ,����  +s����  ,	���F  ,	���F  +s����  +s      D  , ,���p  *���p  *����  *����  *���p  *      D  , ,����  +s����  ,	����  ,	����  +s����  +s      D  , ,��̘  ,���̘  -q���.  -q���.  ,���̘  ,�      D  , ,����  *����  *����  *����  *����  *      D  , ,���X  +s���X  ,	����  ,	����  +s���X  +s      D  , ,���(  *���(  *���ľ  *���ľ  *���(  *      D  , ,����  ,�����  -q���~  -q���~  ,�����  ,�      D  , ,����  ,�����  -q���V  -q���V  ,�����  ,�      D  , ,���   *���   *���Ζ  *���Ζ  *���   *      D  , ,����  +s����  ,	���V  ,	���V  +s����  +s      D  , ,����  *����  *���ǎ  *���ǎ  *����  *      D  , ,����  *����  *����~  *����~  *����  *      D  , ,���   ,����   -q��Ζ  -q��Ζ  ,����   ,�      D  , ,���0  *���0  *�����  *�����  *���0  *      D  , ,���(  +s���(  ,	��ľ  ,	��ľ  +s���(  +s      D  , ,���8  *���8  *�����  *�����  *���8  *      D  , ,����  ,�����  -q���  -q���  ,�����  ,�      D  , ,���p  +s���p  ,	���  ,	���  +s���p  +s      D  , ,���  +s���  ,	����  ,	����  +s���  +s      D  , ,���P  *���P  *�����  *�����  *���P  *      D  , ,��Ő  +s��Ő  ,	���&  ,	���&  +s��Ő  +s      D  , ,���H  +s���H  ,	����  ,	����  +s���H  +s      D  , ,����  ,�����  -q���^  -q���^  ,�����  ,�      D  , ,���H  ,����H  -q����  -q����  ,����H  ,�      D  , ,���h  ,����h  -q����  -q����  ,����h  ,�      D  , ,���   ,����   -q����  -q����  ,����   ,�      D  , ,����  +s����  ,	��ǎ  ,	��ǎ  +s����  +s      D  , ,����  +s����  ,	���~  ,	���~  +s����  +s      D  , ,���P  ,����P  -q����  -q����  ,����P  ,�      D  , ,����  +s����  ,	���  ,	���  +s����  +s      D  , ,���`  +s���`  ,	����  ,	����  +s���`  +s      D  , ,��̘  *��̘  *����.  *����.  *��̘  *      D  , ,���  ,����  -q��՞  -q��՞  ,����  ,�      D  , ,����  ,�����  -q���f  -q���f  ,�����  ,�      D  , ,���(  ,����(  -q��ľ  -q��ľ  ,����(  ,�      D  , ,���  ,����  -q����  -q����  ,����  ,�      D  , ,����  ,�����  -q����  -q����  ,�����  ,�      D  , ,����  +s����  ,	���^  ,	���^  +s����  +s      D  , ,����  *����  *����N  *����N  *����  *      D  , ,����  +s����  ,	���N  ,	���N  +s����  +s      D  , ,���`  *���`  *�����  *�����  *���`  *      D  , ,��Ӡ  +s��Ӡ  ,	���6  ,	���6  +s��Ӡ  +s      D  , ,����  ,�����  -q���F  -q���F  ,�����  ,�      D  , ,���H  *���H  *�����  *�����  *���H  *      D  , ,��Ő  *��Ő  *����&  *����&  *��Ő  *      D  , ,���0  +s���0  ,	����  ,	����  +s���0  +s      D  , ,���   *���   *�����  *�����  *���   *      D  , ,����  +s����  ,	���f  ,	���f  +s����  +s      D  , ,���  *���  *���՞  *���՞  *���  *      D  , ,���8  ,����8  -q����  -q����  ,����8  ,�      D  , ,��Ő  ,���Ő  -q���&  -q���&  ,���Ő  ,�      D  , ,����  *����  *����f  *����f  *����  *      D  , ,���p  ,����p  -q���  -q���  ,����p  ,�      D  , ,��̘  +s��̘  ,	���.  ,	���.  +s��̘  +s      D  , ,����  *����  *����  *����  *����  *      D  , ,����  *����  *����V  *����V  *����  *      D  , ,���8  +s���8  ,	����  ,	����  +s���8  +s      D  , ,����  ,�����  -q���N  -q���N  ,�����  ,�      D  , ,��Ӡ  *��Ӡ  *����6  *����6  *��Ӡ  *      D  , ,����  *����  *����F  *����F  *����  *      D  , ,����  *����  *����^  *����^  *����  *      D  , ,���   +s���   ,	��Ζ  ,	��Ζ  +s���   +s      D  , ,����  *����  *�����  *�����  *����  *      D  , ,���h  *���h  *�����  *�����  *���h  *      D  , ,���`  ,����`  -q����  -q����  ,����`  ,�      D  , ,��Ӡ  ,���Ӡ  -q���6  -q���6  ,���Ӡ  ,�      D  , ,����  ,�����  -q��ǎ  -q��ǎ  ,�����  ,�      D  , ,���X  ,����X  -q����  -q����  ,����X  ,�      D  , ,���  +s���  ,	��՞  ,	��՞  +s���  +s      D  , ,���h  +s���h  ,	����  ,	����  +s���h  +s      D  , ,���X  *���X  *�����  *�����  *���X  *      D  , ,���P  +s���P  ,	����  ,	����  +s���P  +s      D  , ,�������G�����������s�������s���G�������G      D  , ,���k�������k���k������k����������k����      D  , ,���������������k���s���k���s������������      D  , ,���k���G���k�����������������G���k���G      E   ,����������   2����   2���������������      E   ,����  )�����  -�  N�  -�  N�  )�����  )�      E   ,����������   2����   2���������������      E   ,����  )�����  -�  N�  -�  N�  )�����  )�      E     ���e��� VSS       E     ���[  +� VDD       E       N  +� VDD       E        -  +� VDD       E       -�  +� VDD       E     ��ؠ  +� VDD      � 
   % 0� 
   % 0 dac_8bit 
  res_poly$3     ;[   
  res_poly$3     B   
  res_poly$4   �  1)   
  res_poly$3     E   
  res_poly$3     &�   
  res_poly$3   �  	�   
  res_poly$4   �  �   
  res_poly$4   �  
   
  res_poly$4   �  :�   
  res_poly$3   �  Xz   
  res_poly$4   �  NH   
  res_poly$3   	  N�   
  res_poly$4   �  D�   
  res_poly$4   �  W�   
  res_poly$3   �  	�   
  res_poly$3   	  �   
  res_poly$4   �  't      D   ,  �  
�  �  s  h  s  h  
�  �  
�      D   ,  
�  �  
�  (  h  (  h  �  
�  �      D   ,  �  V  �  &�  h  &�  h  V  �  V      D   ,   �  (   �  0�  h  0�  h  (   �  (      D   ,   �  1�   �  :G  h  :G  h  1�   �  1�      D   ,  �  ;u  �  C�  h  C�  h  ;u  �  ;u      D   ,  
�  E*  
�  M�  h  M�  h  E*  
�  E*      D   ,  �  N�  �  Wf  h  Wf  h  N�  �  N�      D   ,   �  <o   �  D�  �  D�  �  <o   �  <o      D   ,  U   �  U  �  �  �  �   �  U   �      D   ,  U  X�  U  `�  �  `�  �  X�  U  X�      D   ,  �   �  �  �  |  �  |   �  �   �      D   ,  
�  
A  
�  y  �  y  �  
A  
�  
A      D   ,  �  �  �  .  �  .  �  �  �  �      D   ,   �  �   �  %�  �  %�  �  �   �  �      D   ,   �  <o   �  D�  �  D�  �  <o   �  <o      D   ,  �  F$  �  N\  �  N\  �  F$  �  F$      D   ,  
�  O�  
�  X  �  X  �  O�  
�  O�      D   ,  �  Y�  �  a�  |  a�  |  Y�  �  Y�      D   ,  �  N�  �  Wf  h  Wf  h  N�  �  N�      D       ;  O� OUT       D       N  S7 OUT       D       	  V� OUT       D         F� DAC5      D         JO DAC5      D         M� DAC5      D         Pn DAC6      D       �  a6 DAC7      D       
�  W� DAC6      D         S� DAC6      D       �  Z' DAC7      D       �  ]� DAC7      D       `  V� OUT       D       [  Sw OUT       D       `  O� OUT       D         D DAC4      D         @� DAC4      D         = DAC4      D          %a DAC3      D       %  !� DAC3      D         I DAC3      D         . DAC2      D         � DAC2      D         � DAC2      D         l DAC1      D         � DAC1      D         
� DAC1      D         � DAC0      D       �  0 DAC0      D       �  * DAC0      D  , ,  �  |  �    @    @  |  �  |      D  , ,  �    �  �  @  �  @    �        D  , ,  �  �  �  B  @  B  @  �  �  �      D  , ,  �  D  �  �  @  �  @  D  �  D      D  , ,  �   �  �  r  @  r  @   �  �   �      D  , ,  �  ^�  �  _  @  _  @  ^�  �  ^�      D  , ,  �  ]  �  ]�  @  ]�  @  ]  �  ]      D  , ,  �  [�  �  \I  @  \I  @  [�  �  [�      D  , ,  �  ZK  �  Z�  @  Z�  @  ZK  �  ZK      D  , ,  �  X�  �  Yy  @  Yy  @  X�  �  X�      D  , ,  �  �  �  {  @  {  @  �  �  �      D  , ,  �  _�  �  `�  @  `�  @  _�  �  _�      E   ,  U   �  U  �  �  �  �   �  U   �      E   ,  U  X�  U  `�  �  `�  �  X�  U  X�      E   ,  U   �  U  �  �  �  �   �  U   �      E   ,  U  X�  U  `�  �  `�  �  X�  U  X�      E       �  `J VDD       E       �  \� VDD       E       �  Y+ VDD       E       �  � VSS       E       �  ! VSS       E       �  , VSS      � 
   % 0� 
   % 0 
driver 
  sky130_fd_sc_hd__buf_16   ?� �   
  sky130_fd_sc_hd__buf_8  *
 �   
  sky130_fd_sc_hd__buf_1  $� �      D   , #� � #� H &c H &c � #� �      D   , e� y e� ! f� ! f� y e� y      C   , )� 0 )� � *� � *� 0 )� 0      C   , ;� 0 ;� � ?� � ?� 0 ;� 0      C   , #� � #� H % H % � #� �      C  , , e� H e� � f� � f� H e� H      C  , , d H d � d� � d� H d H      C  , , e� � e� R f� R f� � e� �      C  , , %� @ %� � &* � &* @ %� @      C  , , d � d R d� R d� � d �      C  , , #� A #� � $� � $� A #� A      C  , , e� � e� � f� � f� � e� �      C  , , e� G e� � f� � f� G e� G      C  , , e� � e� S f� S f� � e� �      C  , , e� Y e�  f�  f� Y e� Y      C  , , e� � e� A f� A f� � e� �      D   , #� � #� H &c H &c � #� �      D   , e� � e�  f�  f� � e� �      D      % � IN      D      fM � OUT       D      fC � OUT       D      fG M OUT       D  , , %A R %A � %� � %� R %A R      D  , , ' R ' � '� � '� R ' R      D  , , *� R *� � +; � +; R *� R      D  , , ,q R ,q � - � - R ,q R      D  , , .= R .= � .� � .� R .= R      D  , , 0	 R 0	 � 0� � 0� R 0	 R      D  , , 1� R 1� � 2k � 2k R 1� R      D  , , (� R (� � )o � )o R (� R      D  , , 3� R 3� � 47 � 47 R 3� R      D  , , 5m R 5m � 6 � 6 R 5m R      D  , , 9 R 9 � 9� � 9� R 9 R      D  , , :� R :� � ;g � ;g R :� R      D  , , <� R <� � =3 � =3 R <� R      D  , , >i R >i � >� � >� R >i R      D  , , @5 R @5 � @� � @� R @5 R      D  , , 79 R 79 � 7� � 7� R 79 R      D  , , B R B � B� � B� R B R      D  , , C� R C� � Dc � Dc R C� R      D  , , Ge R Ge � G� � G� R Ge R      D  , , I1 R I1 � I� � I� R I1 R      D  , , J� R J� � K� � K� R J� R      D  , , L� R L� � M_ � M_ R L� R      D  , , N� R N� � O+ � O+ R N� R      D  , , E� R E� � F/ � F/ R E� R      D  , , Pa R Pa � P� � P� R Pa R      D  , , R- R R- � R� � R� R R- R      D  , , U� R U� � V[ � V[ R U� R      D  , , W� R W� � X' � X' R W� R      D  , , Y] R Y] � Y� � Y� R Y] R      D  , , [) R [) � [� � [� R [) R      D  , , \� R \� � ]� � ]� R \� R      D  , , S� R S� � T� � T� R S� R      D  , , ^� R ^� � _W � _W R ^� R      D  , , `� R `� � a# � a# R `� R      D  , , bY R bY � b� � b� R bY R      D  , , d% R d% � d� � d� R d% R      D  , , e� R e� � f� � f� R e� R      D  , , %A � %A H %� H %� � %A �      D  , , ' � ' H '� H '� � ' �      D  , , *� � *� H +; H +; � *� �      D  , , ,q � ,q H - H - � ,q �      D  , , .= � .= H .� H .� � .= �      D  , , 0	 � 0	 H 0� H 0� � 0	 �      D  , , 1� � 1� H 2k H 2k � 1� �      D  , , (� � (� H )o H )o � (� �      D  , , 3� � 3� H 47 H 47 � 3� �      D  , , 5m � 5m H 6 H 6 � 5m �      D  , , 9 � 9 H 9� H 9� � 9 �      D  , , :� � :� H ;g H ;g � :� �      D  , , <� � <� H =3 H =3 � <� �      D  , , >i � >i H >� H >� � >i �      D  , , @5 � @5 H @� H @� � @5 �      D  , , 79 � 79 H 7� H 7� � 79 �      D  , , B � B H B� H B� � B �      D  , , C� � C� H Dc H Dc � C� �      D  , , Ge � Ge H G� H G� � Ge �      D  , , I1 � I1 H I� H I� � I1 �      D  , , J� � J� H K� H K� � J� �      D  , , L� � L� H M_ H M_ � L� �      D  , , N� � N� H O+ H O+ � N� �      D  , , E� � E� H F/ H F/ � E� �      D  , , Pa � Pa H P� H P� � Pa �      D  , , R- � R- H R� H R� � R- �      D  , , U� � U� H V[ H V[ � U� �      D  , , W� � W� H X' H X' � W� �      D  , , Y] � Y] H Y� H Y� � Y] �      D  , , [) � [) H [� H [� � [) �      D  , , \� � \� H ]� H ]� � \� �      D  , , S� � S� H T� H T� � S� �      D  , , ^� � ^� H _W H _W � ^� �      D  , , `� � `� H a# H a# � `� �      D  , , bY � bY H b� H b� � bY �      D  , , d% � d% H d� H d� � d% �      D  , , e� � e� H f� H f� � e� �      E   , $� � $� � g" � g" � $� �      E   , $�  $� � g" � g"  $�       E   , $� � $� � g" � g" � $� �      E   , $�  $� � g" � g"  $�       E      %b � VSS       E      fd  VSS       E      E�  VSS       E      32  VSS       E      W� , VSS       E      %� � VDD       E      f# � VDD       E      E� � VDD       E      3] � VDD       E      X � VDD      � 
   % 0� 
   % 0 tt_um_template       , � �� � ��  ��  �� � ��         , � �� � �� � �� � �� � ��         ,  ��  �� J �� J ��  ��         , �V �� �V �� �� �� �� �� �V ��         , � �� � �� � �� � �� � ��         , �� �� �� �� �� �� �� �� �� ��         , �� �� �� �� �* �� �* �� �� ��         , �6 �� �6 �� �b �� �b �� �6 ��         , �n �� �n �� Ú �� Ú �� �n ��         , �� �� �� �� �� �� �� �� �� ��         , �� �� �� �� �
 �� �
 �� �� ��         , � �� � �� �B �� �B �� � ��         , �N �� �N �� �z �� �z �� �N ��         , �� �� �� �� �� �� �� �� �� ��         , �� �� �� �� �� �� �� �� �� ��         , v� �� v� �� x" �� x" �� v� ��         , l. �� l. �� mZ �� mZ �� l. ��         , af �� af �� b� �� b� �� af ��         , V� �� V� �� W� �� W� �� V� ��         ,  �V ��  �V ��  �� ��  �� ��  �V ��         ,  �� ��  �� ��  �� ��  �� ��  �� ��         ,  �� ��  �� ��  �� ��  �� ��  �� ��         ,  ~� ��  ~� ��  �* ��  �* ��  ~� ��         ,  t6 ��  t6 ��  ub ��  ub ��  t6 ��         ,  in ��  in ��  j� ��  j� ��  in ��         ,  ^� ��  ^� ��  _� ��  _� ��  ^� ��         ,  S� ��  S� ��  U
 ��  U
 ��  S� ��         ,  �� ��  �� ��  �� ��  �� ��  �� ��         ,  �� ��  �� ��  �� ��  �� ��  �� ��         ,  � ��  � ��  �2 ��  �2 ��  � ��         ,  �> ��  �> ��  �j ��  �j ��  �> ��         ,  �v ��  �v ��  ˢ ��  ˢ ��  �v ��         ,  �� ��  �� ��  �� ��  �� ��  �� ��         ,  �� ��  �� ��  � ��  � ��  �� ��         ,  � ��  � ��  �J ��  �J ��  � ��         , K� �� K� �� M �� M �� K� ��         , A �� A �� B: �� B: �� A ��         , 6F �� 6F �� 7r �� 7r �� 6F ��         , +~ �� +~ �� ,� �� ,� �� +~ ��         ,  � ��  � �� !� �� !� ��  � ��         , � �� � ��  ��  �� � ��         , & �� & �� R �� R �� & ��         ,  ^ ��  ^ �� � �� � ��  ^ ��          ,             �� f� �� f�                      | �� clk           D �� ena           � �� 
rst_n           �� �� ui_in[0]          �$ �� ui_in[1]          �\ �� ui_in[2]          ؔ �� ui_in[3]          �� �� ui_in[4]          � �� ui_in[5]          �< �� ui_in[6]          �t �� ui_in[7]          �� �� uio_in[0]           �� �� uio_in[1]           � �� uio_in[2]           �T �� uio_in[3]           w� �� uio_in[4]           l� �� uio_in[5]           a� �� uio_in[6]           W4 �� uio_in[7]            �� �� uio_oe[0]            �$ �� uio_oe[1]            �\ �� uio_oe[2]            � �� uio_oe[3]            t� �� uio_oe[4]            j �� uio_oe[5]            _< �� uio_oe[6]            Tt �� uio_oe[7]            �, �� uio_out[0]           �d �� uio_out[1]           �� �� uio_out[2]           �� �� uio_out[3]           � �� uio_out[4]           �D �� uio_out[5]           �| �� uio_out[6]           �� �� uio_out[7]          Ll �� uo_out[0]           A� �� uo_out[1]           6� �� uo_out[2]           , �� uo_out[3]           !L �� uo_out[4]           � �� uo_out[5]           � �� uo_out[6]            � �� uo_out[7]      � 
   % 0� 
   % 0 pin_connect     D   ,              �  r  �  r                  D  , ,   n  �   n  b    b    �   n  �      D  , ,   n   n   n           n   n   n      E   ,����    ����  �  w  �  w    ����          F  , ,   U  J   U          J   U  J      F  , ,   U  �   U  �    �    �   U  �      E  , ,   U  �   U  �    �    �   U  �      E  , ,   U  *   U  �    �    *   U  *      G   ,����  �����  �  w  �  w  �����  �      G   ,   #  �   #  
   O  
   O  �   #  �      F   ,����  �����  �  w  �  w  �����  �     � 
   % 0� 
   % 0 tt_um_wulf_8bit_vco  
  dac_8bit �  C�       �� ��   
  inv_strvd  �  B�        �� -   
  
driver    B�        ]� ��   
  inv_strvd  �  BZ         �� �P   
  inv_strvd  �  C�       Z@ �X   
  inv_strvd  �  B�        Y� �   
  inv_strvd  �   �  v�   
  inv_strvd  �   #f ~_   
  inv_strvd  �  BZ         �q U�   
  pin_connect    �� �b   
  pin_connect   � �b   
  pin_connect   J �b   
  pin_connect    �b   
  pin_connect   '� �b   
  pin_connect   2� �b   
  pin_connect   =j �b   
  pin_connect   H2 �b   
  pin_connect   R� �b   
  pin_connect   ]� �b   
  pin_connect   h� �b   
  pin_connect   sR �b   
  pin_connect   ~ �b   
  pin_connect   �� �b   
  pin_connect   �� �b   
  pin_connect   �r �b   
  pin_connect   �: �b   
  pin_connect   � �b   
  pin_connect   �� �b   
  pin_connect   ɒ �b   
  pin_connect   �Z �b   
  pin_connect   �" �b   
  pin_connect   �� �b   
  pin_connect   �� �b   
  pin_connect   �z �b   
  pin_connect   
B �b   
  pin_connect   
 �b   
  pin_connect   � �b   
  pin_connect   *� �b   
  pin_connect   5b �b   
  pin_connect   @* �b   
  pin_connect   J� �b   
  pin_connect   U� �b   
  pin_connect   `� �b   
  pin_connect   kJ �b   
  pin_connect   v �b   
  pin_connect   �� �b   
  pin_connect   �� �b   
  pin_connect   �j �b   
  pin_connect   �2 �b   
  pin_connect   �� �b   
  pin_connect   �� �b   
  pin_connect   �� �b   
  tt_um_template   ��  ��      D   , `� &� `� J� i� J� i� &� `� &�      D   , �G  �G 	� DJ 	� DJ  �G       D   ,  �� ��  �� ��  �T ��  �T ��  �� ��      D   , :� a� :� �a <7 �a <7 a� :� a�      D   , [� �6 [� �b a� �b a� �6 [� �6      D   ,  �� ��  �� �a �a �a �a ��  �� ��      D   , T� �b T� �� \� �� \� �b T� �b      D   , ^D �X ^D �� f| �� f| �X ^D �X      D   , Q� �6 Q� �b W, �b W, �6 Q� �6      D   , eP �6 eP �b l� �b l� �6 eP �6      D   , �j �6 �j �b �S �b �S �6 �j �6      D   , �� �6 �� �b �� �b �� �6 �� �6      D   , g� �N g� �z p1 �z p1 �N g� �N      D   , o �6 o �b w� �b w� �6 o �6      D   , �' �b �' �� �_ �� �_ �b �' �b      D   , �� �l �� �� � �� � �l �� �l      D   , �2 �6 �2 �b � �b � �6 �2 �6      D   , �� �6 �� �b �� �b �� �6 �� �6      D   , �� �� �� �6 � �6 � �� �� ��      D   , �r �� �r �6 �� �6 �� �� �r ��      D   , �� �N �� �z �� �z �� �N �� �N      D   , �' �� �' �6 �S �6 �S �� �' ��      D   , �r �X �r �� �� �� �� �X �r �X      D   , �� �z �� �6 �� �6 �� �z �� �z      D   , o �z o �6 p1 �6 p1 �z o �z      D   , eP �� eP �6 f| �6 f| �� eP ��      D   , [� �� [� �6 \� �6 \� �� [� ��      D   , Q� �� Q� �6 S �6 S �� Q� ��      D   , J� �l J� �� S �� S �l J� �l      D   , 9� �a 9� �� <7 �� <7 �a 9� �a      D   , �� �� �� �b �$ �b �$ �� �� ��      D   , �$ �� �$ �0 �% �0 �% �� �$ ��      D   , "� a� "� i� :� i� :� a� "� a�      D   , 5L M� 5L a� :� a� :� M� 5L M�      D   , ]� J� ]� S~ i� S~ i� J� ]� J�      D   , U: J� U: w� ]� w� ]� J� U: J�      D   , r: h� r: p� �� p� �� h� r: h�      D   ,  �T |T  �T ��  �� ��  �� |T  �T |T      D   ,  �A ��  �A �a  �� �a  �� ��  �A ��      D   , }� t� }� �� �a �� �a t� }� t�      D   ,  �? E$  �? x[  �7 x[  �7 E$  �? E$      D   ,  �u �  �u � � � � �  �u �      D   , �� � �� :� �� :� �� � �� �      D   ,  �|  �  �|  �� �G  �� �G  �  �|  �      D   ,  ��  �  ��  ��  �|  ��  �|  �  ��  �      D   ,  �T  ��  �T %  �| %  �|  ��  �T  ��      D   ,  �T %  �T ��  �� ��  �� %  �T %      D   ,  �� �*  �� ��  �T ��  �T �*  �� �*      D   , �G  � �G  ��  ��  � �G  �      D   ,  �� �)  �� �!  �� �!  �� �)  �� �)      D   , 
� � 
�  �  � � 
� �      D   , DJ &� DJ / `� / `� &� DJ &�      D   , DJ  DJ &� L� &� L�  DJ       D   , D� 3 D� �� L� �� L� 3 D� 3      E   , ��  �� �� N� K� N� K�  �� ��  ��      E   ,  ��  ��  �� J�  � J�  �  ��  ��  ��      E   ,  �y \+  �y �B B �B B \+  �y \+      E   ,  � ��  � A #� A #� ��  � ��      E   , �� b� �� �� #� �� #� b� �� b�      E   , R� �B R� �9 �a �9 �a �B R� �B      E   ,  �� \+  �� ��  �y ��  �y \+  �� \+      E   ,  � �  � ��  �� ��  �� �  � �      E   , � U � z+ C� z+ C� U � U      E   , A" z+ A" �� C� �� C� z+ A" z+      E   , #� b� #� �� K� �� K� b� #� b�      E   , 8d �� 8d U K� U K� �� 8d ��      E   ,  �� J�  �� \+  �x \+  �x J�  �� J�      E   ,  �W A  �W H� y� H� y� A  �W A      E   ,  �W ��  �W A  � A  � ��  �W ��      E   ,  �W ��  �W ��  �� ��  �� ��  �W ��      E   , y� A y� \+ B \+ B A y� A      E   , �� =� �� N� �� N� �� =� �� =�      E   , C� U C� t� K� t� K� U C� U      E   ,  �  ��  � � < � <  ��  �  ��      E   , �9 t� �9 �� � �� � t� �9 t�      E   , K� |@ K� }� T+ }� T+ |@ K� |@      E   , <  �� < )� �� )� ��  �� <  ��      E   , < =� < �� �� �� �� =� < =�      E   , [ t� [ �� �9 �� �9 t� [ t�      E   , A" �� A" �B �9 �B �9 �� A" ��      E   , K�  �� K� t� � t� �  �� K�  ��      E   , B U B �B � �B � U B U      E   , � �P � �B A" �B A" �P � �P      F  , , � 3� � 4� 	� 4� 	� 3� � 3�      F  , , � 3� � 4� [ 4� [ 3� � 3�      F  , ,  3�  4� � 4� � 3�  3�      F  , , 
s 3� 
s 4� ; 4� ; 3� 
s 3�      F  , , � �& � �� 	� �� 	� �& � �&      F  , ,  �&  �� � �� � �&  �&      F  , , 
s �& 
s �� ; �� ; �& 
s �&      F  , , � �& � �� [ �� [ �& � �&      F  , , � �6 � �� [ �� [ �6 � �6      F  , , 
s �& 
s �� ; �� ; �& 
s �&      F  , , � �� � �� [ �� [ �� � ��      F  , , 
s �� 
s �~ ; �~ ; �� 
s ��      F  , , � �V � � [ � [ �V � �V      F  , , � �� � �� [ �� [ �� � ��      F  , , � �v � �> [ �> [ �v � �v      F  , , � � � �� [ �� [ � � �      F  , , � �� � �^ [ �^ [ �� � ��      F  , , 
s �V 
s � ; � ; �V 
s �V      F  , , � �& � �� [ �� [ �& � �&      F  , , � �� � �~ 	� �~ 	� �� � ��      F  , , � �� � �~ [ �~ [ �� � ��      F  , , � �F � � 	� � 	� �F � �F      F  , , � �� � �� 	� �� 	� �� � ��      F  , , � �f � �. 	� �. 	� �f � �f      F  , , � �� � �� 	� �� 	� �� � ��      F  , , � �� � �N 	� �N 	� �� � ��      F  , , � �� � �� [ �� [ �� � ��      F  , , � � � �� 	� �� 	� � � �      F  , ,  ��  �~ � �~ � ��  ��      F  , , � �� � �n 	� �n 	� �� � ��      F  , ,  �F  � � � � �F  �F      F  , , � �6 � �� 	� �� 	� �6 � �6      F  , ,  ��  �� � �� � ��  ��      F  , , � �� � �� 	� �� 	� �� � ��      F  , ,  �f  �. � �. � �f  �f      F  , , 
s �v 
s �> ; �> ; �v 
s �v      F  , , � �V � � 	� � 	� �V � �V      F  , ,  ��  �� � �� � ��  ��      F  , , � �� � �� 	� �� 	� �� � ��      F  , ,  ��  �N � �N � ��  ��      F  , , � �v � �> 	� �> 	� �v � �v      F  , ,  �  �� � �� � �  �      F  , , � � � �� 	� �� 	� � � �      F  , ,  ��  �n � �n � ��  ��      F  , , � �� � �^ 	� �^ 	� �� � ��      F  , ,  �6  �� � �� � �6  �6      F  , , � �& � �� 	� �� 	� �& � �&      F  , ,  ��  �� � �� � ��  ��      F  , , � �� � �~ 	� �~ 	� �� � ��      F  , ,  �V  � � � � �V  �V      F  , ,  ��  �� � �� � ��  ��      F  , ,  �v  �> � �> � �v  �v      F  , ,  �  �� � �� � �  �      F  , ,  ��  �^ � �^ � ��  ��      F  , ,  �&  �� � �� � �&  �&      F  , ,  ��  �~ � �~ � ��  ��      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , , 
s �� 
s �~ ; �~ ; �� 
s ��      F  , , 
s �F 
s � ; � ; �F 
s �F      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , , 
s �f 
s �. ; �. ; �f 
s �f      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , , 
s �� 
s �N ; �N ; �� 
s ��      F  , , � �� � �N [ �N [ �� � ��      F  , , 
s � 
s �� ; �� ; � 
s �      F  , , � �� � �~ [ �~ [ �� � ��      F  , , 
s �� 
s �n ; �n ; �� 
s ��      F  , , � �F � � [ � [ �F � �F      F  , , 
s �6 
s �� ; �� ; �6 
s �6      F  , , � �� � �� [ �� [ �� � ��      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , , � �f � �. [ �. [ �f � �f      F  , , � � � �� [ �� [ � � �      F  , , 
s � 
s �� ; �� ; � 
s �      F  , , � �� � �n [ �n [ �� � ��      F  , , 
s �� 
s �^ ; �^ ; �� 
s ��      F  , , 
s p� 
s q� ; q� ; p� 
s p�      F  , ,  oF  p � p � oF  oF      F  , , � ~� � � [ � [ ~� � ~�      F  , , � z6 � z� 	� z� 	� z6 � z6      F  , ,  j�  k^ � k^ � j�  j�      F  , ,  p�  q� � q� � p�  p�      F  , , 
s rf 
s s. ; s. ; rf 
s rf      F  , , � {� � |� 	� |� 	� {� � {�      F  , , � �v � �> [ �> [ �v � �v      F  , ,  rf  s. � s. � rf  rf      F  , , � s� � t� 	� t� 	� s� � s�      F  , , � }V � ~ 	� ~ 	� }V � }V      F  , , 
s s� 
s t� ; t� ; s� 
s s�      F  , ,  s�  t� � t� � s�  s�      F  , , � ~� � � 	� � 	� ~� � ~�      F  , , � � � �� [ �� [ � � �      F  , ,  u�  vN � vN � u�  u�      F  , , � �v � �> 	� �> 	� �v � �v      F  , , 
s u� 
s vN ; vN ; u� 
s u�      F  , ,  w  w� � w� � w  w      F  , , � � � �� 	� �� 	� � � �      F  , , � oF � p 	� p 	� oF � oF      F  , ,  x�  yn � yn � x�  x�      F  , , � �� � �^ 	� �^ 	� �� � ��      F  , ,  l&  l� � l� � l&  l&      F  , , 
s w 
s w� ; w� ; w 
s w      F  , ,  z6  z� � z� � z6  z6      F  , , � j� � k^ 	� k^ 	� j� � j�      F  , , 
s x� 
s yn ; yn ; x� 
s x�      F  , ,  {�  |� � |� � {�  {�      F  , , � j� � k^ [ k^ [ j� � j�      F  , , � �� � �^ [ �^ [ �� � ��      F  , ,  }V  ~ � ~ � }V  }V      F  , , � l& � l� [ l� [ l& � l&      F  , ,  ~�  � � � � ~�  ~�      F  , , 
s z6 
s z� ; z� ; z6 
s z6      F  , ,  �v  �> � �> � �v  �v      F  , , � m� � n~ [ n~ [ m� � m�      F  , ,  �  �� � �� � �  �      F  , , � rf � s. 	� s. 	� rf � rf      F  , ,  ��  �^ � �^ � ��  ��      F  , , 
s {� 
s |� ; |� ; {� 
s {�      F  , , � oF � p [ p [ oF � oF      F  , , � l& � l� 	� l� 	� l& � l&      F  , , 
s }V 
s ~ ; ~ ; }V 
s }V      F  , , � p� � q� [ q� [ p� � p�      F  , , 
s ~� 
s � ; � ; ~� 
s ~�      F  , , � rf � s. [ s. [ rf � rf      F  , , � s� � t� [ t� [ s� � s�      F  , , 
s �v 
s �> ; �> ; �v 
s �v      F  , , � u� � vN [ vN [ u� � u�      F  , , 
s � 
s �� ; �� ; � 
s �      F  , , � w � w� [ w� [ w � w      F  , , 
s �� 
s �^ ; �^ ; �� 
s ��      F  , , 
s j� 
s k^ ; k^ ; j� 
s j�      F  , , � x� � yn [ yn [ x� � x�      F  , , � w � w� 	� w� 	� w � w      F  , , 
s l& 
s l� ; l� ; l& 
s l&      F  , , � u� � vN 	� vN 	� u� � u�      F  , , � z6 � z� [ z� [ z6 � z6      F  , , 
s m� 
s n~ ; n~ ; m� 
s m�      F  , , � {� � |� [ |� [ {� � {�      F  , , � p� � q� 	� q� 	� p� � p�      F  , , 
s oF 
s p ; p ; oF 
s oF      F  , , � }V � ~ [ ~ [ }V � }V      F  , ,  m�  n~ � n~ � m�  m�      F  , , � m� � n~ 	� n~ 	� m� � m�      F  , , � x� � yn 	� yn 	� x� � x�      F  , , � Nv � O> 	� O> 	� Nv � Nv      F  , , 
s Nv 
s O> ; O> ; Nv 
s Nv      F  , , � Nv � O> [ O> [ Nv � Nv      F  , ,  Nv  O> � O> � Nv  Nv      F  , , � W� � X� 	� X� 	� W� � W�      F  , , 
s _� 
s `n ; `n ; _� 
s _�      F  , , � e� � f� 	� f� 	� e� � e�      F  , , 
s a6 
s a� ; a� ; a6 
s a6      F  , ,  _�  `n � `n � _�  _�      F  , ,  b�  c� � c� � b�  b�      F  , , 
s b� 
s c� ; c� ; b� 
s b�      F  , , � Yf � Z. 	� Z. 	� Yf � Yf      F  , , � P � P� [ P� [ P � P      F  , ,  \�  ]N � ]N � \�  \�      F  , , 
s dV 
s e ; e ; dV 
s dV      F  , , � Q� � R^ [ R^ [ Q� � Q�      F  , , 
s e� 
s f� ; f� ; e� 
s e�      F  , , � S& � S� [ S� [ S& � S&      F  , , � Z� � [� 	� [� 	� Z� � Z�      F  , , � T� � U~ [ U~ [ T� � T�      F  , , 
s gv 
s h> ; h> ; gv 
s gv      F  , , � gv � h> 	� h> 	� gv � gv      F  , , � VF � W [ W [ VF � VF      F  , ,  T�  U~ � U~ � T�  T�      F  , , 
s i 
s i� ; i� ; i 
s i      F  , ,  ^  ^� � ^� � ^  ^      F  , , � W� � X� [ X� [ W� � W�      F  , , � \� � ]N 	� ]N 	� \� � \�      F  , ,  P  P� � P� � P  P      F  , , � Yf � Z. [ Z. [ Yf � Yf      F  , ,  Q�  R^ � R^ � Q�  Q�      F  , , � ^ � ^� 	� ^� 	� ^ � ^      F  , , � Z� � [� [ [� [ Z� � Z�      F  , , � i � i� 	� i� 	� i � i      F  , , � \� � ]N [ ]N [ \� � \�      F  , ,  S&  S� � S� � S&  S&      F  , , 
s \� 
s ]N ; ]N ; \� 
s \�      F  , ,  Z�  [� � [� � Z�  Z�      F  , ,  e�  f� � f� � e�  e�      F  , , 
s ^ 
s ^� ; ^� ; ^ 
s ^      F  , , 
s Q� 
s R^ ; R^ ; Q� 
s Q�      F  , , � b� � c� 	� c� 	� b� � b�      F  , , � Q� � R^ 	� R^ 	� Q� � Q�      F  , , 
s S& 
s S� ; S� ; S& 
s S&      F  , , � e� � f� [ f� [ e� � e�      F  , ,  W�  X� � X� � W�  W�      F  , , 
s T� 
s U~ ; U~ ; T� 
s T�      F  , , � S& � S� 	� S� 	� S& � S&      F  , , � gv � h> [ h> [ gv � gv      F  , , 
s VF 
s W ; W ; VF 
s VF      F  , ,  gv  h> � h> � gv  gv      F  , , � T� � U~ 	� U~ 	� T� � T�      F  , , 
s W� 
s X� ; X� ; W� 
s W�      F  , , � i � i� [ i� [ i � i      F  , ,  Yf  Z. � Z. � Yf  Yf      F  , , 
s Yf 
s Z. ; Z. ; Yf 
s Yf      F  , , � dV � e 	� e 	� dV � dV      F  , , � VF � W 	� W 	� VF � VF      F  , , 
s Z� 
s [� ; [� ; Z� 
s Z�      F  , ,  i  i� � i� � i  i      F  , , � P � P� 	� P� 	� P � P      F  , , 
s P 
s P� ; P� ; P 
s P      F  , ,  a6  a� � a� � a6  a6      F  , , � dV � e [ e [ dV � dV      F  , , � _� � `n [ `n [ _� � _�      F  , ,  dV  e � e � dV  dV      F  , , � a6 � a� 	� a� 	� a6 � a6      F  , , � ^ � ^� [ ^� [ ^ � ^      F  , , � a6 � a� [ a� [ a6 � a6      F  , ,  VF  W � W � VF  VF      F  , , � _� � `n 	� `n 	� _� � _�      F  , , � b� � c� [ c� [ b� � b�      F  , , � =F � > 	� > 	� =F � =F      F  , , 
s L� 
s M� ; M� ; L� 
s L�      F  , , � 8� � 9^ [ 9^ [ 8� � 8�      F  , , � ;� � <~ 	� <~ 	� ;� � ;�      F  , , � L� � M� [ M� [ L� � L�      F  , , 
s I� 
s J� ; J� ; I� 
s I�      F  , ,  @f  A. � A. � @f  @f      F  , ,  =F  > � > � =F  =F      F  , ,  8�  9^ � 9^ � 8�  8�      F  , , � >� � ?� [ ?� [ >� � >�      F  , ,  KV  L � L � KV  KV      F  , , � I� � J� [ J� [ I� � I�      F  , , � >� � ?� 	� ?� 	� >� � >�      F  , ,  >�  ?� � ?� � >�  >�      F  , , � F� � Gn 	� Gn 	� F� � F�      F  , , � =F � > [ > [ =F � =F      F  , ,  A�  B� � B� � A�  A�      F  , ,  ;�  <~ � <~ � ;�  ;�      F  , , � 5v � 6> [ 6> [ 5v � 5v      F  , ,  5v  6> � 6> � 5v  5v      F  , , � @f � A. 	� A. 	� @f � @f      F  , ,  C�  DN � DN � C�  C�      F  , , � L� � M� 	� M� 	� L� � L�      F  , , 
s 5v 
s 6> ; 6> ; 5v 
s 5v      F  , , � ;� � <~ [ <~ [ ;� � ;�      F  , , 
s C� 
s DN ; DN ; C� 
s C�      F  , ,  L�  M� � M� � L�  L�      F  , ,  E  E� � E� � E  E      F  , , � A� � B� 	� B� 	� A� � A�      F  , , � @f � A. [ A. [ @f � @f      F  , , 
s >� 
s ?� ; ?� ; >� 
s >�      F  , , � H6 � H� 	� H� 	� H6 � H6      F  , , 
s E 
s E� ; E� ; E 
s E      F  , , 
s H6 
s H� ; H� ; H6 
s H6      F  , , � 5v � 6> 	� 6> 	� 5v � 5v      F  , , � A� � B� [ B� [ A� � A�      F  , ,  F�  Gn � Gn � F�  F�      F  , , 
s :& 
s :� ; :� ; :& 
s :&      F  , , � 7 � 7� [ 7� [ 7 � 7      F  , , � C� � DN 	� DN 	� C� � C�      F  , , � C� � DN [ DN [ C� � C�      F  , , � 7 � 7� 	� 7� 	� 7 � 7      F  , , 
s 7 
s 7� ; 7� ; 7 
s 7      F  , ,  7  7� � 7� � 7  7      F  , , � E � E� [ E� [ E � E      F  , , 
s ;� 
s <~ ; <~ ; ;� 
s ;�      F  , ,  H6  H� � H� � H6  H6      F  , , � 8� � 9^ 	� 9^ 	� 8� � 8�      F  , , � F� � Gn [ Gn [ F� � F�      F  , , � :& � :� [ :� [ :& � :&      F  , ,  :&  :� � :� � :&  :&      F  , , � E � E� 	� E� 	� E � E      F  , , � :& � :� 	� :� 	� :& � :&      F  , , � H6 � H� [ H� [ H6 � H6      F  , , � KV � L 	� L 	� KV � KV      F  , , � I� � J� 	� J� 	� I� � I�      F  , , 
s 8� 
s 9^ ; 9^ ; 8� 
s 8�      F  , , 
s =F 
s > ; > ; =F 
s =F      F  , , � KV � L [ L [ KV � KV      F  , , 
s KV 
s L ; L ; KV 
s KV      F  , , 
s F� 
s Gn ; Gn ; F� 
s F�      F  , , 
s @f 
s A. ; A. ; @f 
s @f      F  , , 
s A� 
s B� ; B� ; A� 
s A�      F  , ,  I�  J� � J� � I�  I�      F  , ,  �6  �� � �� � �6  �6      F  , , 
s �6 
s �� ; �� ; �6 
s �6      F  , , � �6 � �� [ �� [ �6 � �6      F  , , � �6 � �� 	� �� 	� �6 � �6      F  , , 
s  
s � ; � ;  
s       F  , , � "� � #~ [ #~ [ "� � "�      F  , ,  "�  #~ � #~ � "�  "�      F  , , � $F � % [ % [ $F � $F      F  , ,  $F  % � % � $F  $F      F  , , � %� � &� [ &� [ %� � %�      F  , ,  %�  &� � &� � %�  %�      F  , , 
s � 
s  ^ ;  ^ ; � 
s �      F  , , � 'f � (. [ (. [ 'f � 'f      F  , ,  'f  (. � (. � 'f  'f      F  , , 
s !& 
s !� ; !� ; !& 
s !&      F  , , � � � � 	� � 	� � � �      F  , , � (� � )� [ )� [ (� � (�      F  , ,  (�  )� � )� � (�  (�      F  , , � *� � +N [ +N [ *� � *�      F  , ,  *�  +N � +N � *�  *�      F  , , 
s "� 
s #~ ; #~ ; "� 
s "�      F  , , � , � ,� [ ,� [ , � ,      F  , ,  ,  ,� � ,� � ,  ,      F  , , � %� � &� 	� &� 	� %� � %�      F  , , � -� � .n [ .n [ -� � -�      F  , ,  -�  .n � .n � -�  -�      F  , , 
s $F 
s % ; % ; $F 
s $F      F  , , � /6 � /� [ /� [ /6 � /6      F  , ,  /6  /� � /� � /6  /6      F  , , � !& � !� 	� !� 	� !& � !&      F  , , � v � > 	� > 	� v � v      F  , , 
s %� 
s &� ; &� ; %� 
s %�      F  , , � 0� � 1� [ 1� [ 0� � 0�      F  , ,  0�  1� � 1� � 0�  0�      F  , , � 2V � 3 [ 3 [ 2V � 2V      F  , ,  2V  3 � 3 � 2V  2V      F  , , � $F � % 	� % 	� $F � $F      F  , , 
s 'f 
s (. ; (. ; 'f 
s 'f      F  , , 
s (� 
s )� ; )� ; (� 
s (�      F  , , 
s *� 
s +N ; +N ; *� 
s *�      F  , , �  � � 	� � 	�  �       F  , , � !& � !� [ !� [ !& � !&      F  , ,  !&  !� � !� � !&  !&      F  , , 
s 2V 
s 3 ; 3 ; 2V 
s 2V      F  , , � (� � )� 	� )� 	� (� � (�      F  , , � *� � +N 	� +N 	� *� � *�      F  , , 
s -� 
s .n ; .n ; -� 
s -�      F  , , � , � ,� 	� ,� 	� , � ,      F  , , � 'f � (. 	� (. 	� 'f � 'f      F  , , � "� � #~ 	� #~ 	� "� � "�      F  , ,  V   �  � V  V      F  , , � -� � .n 	� .n 	� -� � -�      F  , , 
s V 
s  ;  ; V 
s V      F  , , � /6 � /� 	� /� 	� /6 � /6      F  , , 
s /6 
s /� ; /� ; /6 
s /6      F  , , � 0� � 1� 	� 1� 	� 0� � 0�      F  , , � V �  [  [ V � V      F  , ,  �  � � � � �  �      F  , , 
s � 
s � ; � ; � 
s �      F  , , � � � � [ � [ � � �      F  , , � 2V � 3 	� 3 	� 2V � 2V      F  , , � v � > [ > [ v � v      F  , , � V �  	�  	� V � V      F  , , �  � � [ � [  �       F  , ,    � � � �         F  , , 
s 0� 
s 1� ; 1� ; 0� 
s 0�      F  , ,  v  > � > � v  v      F  , , 
s v 
s > ; > ; v 
s v      F  , , � � �  ^ [  ^ [ � � �      F  , ,  �   ^ �  ^ � �  �      F  , , 
s , 
s ,� ; ,� ; , 
s ,      F  , , � � �  ^ 	�  ^ 	� � � �      F  , , � � � � [ � [ � � �      F  , , 
s � 
s N ; N ; � 
s �      F  , ,   V   �  �  V   V      F  , ,  �  � � � � �  �      F  , , 
s  V 
s  ;  ;  V 
s  V      F  , , � � � � 	� � 	� � � �      F  , , 
s � 
s � ; � ; � 
s �      F  , ,  �  � � � � �  �      F  , , 
s � 
s � ; � ; � 
s �      F  , ,    � � � �         F  , , 
s 6 
s � ; � ; 6 
s 6      F  , ,  �  � � � � �  �      F  , , � � � N [ N [ � � �      F  , , 
s � 
s � ; � ; � 
s �      F  , , � 	� � 
~ [ 
~ [ 	� � 	�      F  , , 
s  
s � ; � ;  
s       F  , , � & � � 	� � 	� & � &      F  , , � � � ^ 	� ^ 	� � � �      F  , , � F �  	�  	� F � F      F  , ,  v  > � > � v  v      F  , , 
s v 
s > ; > ; v 
s v      F  , , �  � � [ � [  �       F  , , � 	� � 
~ 	� 
~ 	� 	� � 	�      F  , , � � � � [ � [ � � �      F  , , � � � N 	� N 	� � � �      F  , , � v � > 	� > 	� v � v      F  , , � � � n 	� n 	� � � �      F  , , 
s  
s � ; � ;  
s       F  , , 
s � 
s � ; � ; � 
s �      F  , , 
s � 
s n ; n ; � 
s �      F  , ,  f  . � . � f  f      F  , , �  V �  	�  	�  V �  V      F  , , 
s & 
s � ; � ; & 
s &      F  , , � � � n [ n [ � � �      F  , ,  6  � � � � 6  6      F  , ,  	�  
~ � 
~ � 	�  	�      F  , , � & � � [ � [ & � &      F  , , � 6 � � 	� � 	� 6 � 6      F  , , �  � � 	� � 	�  �       F  , , � �� � �� 	� �� 	� �� � ��      F  , ,  �  n � n � �  �      F  , , 
s 	� 
s 
~ ; 
~ ; 	� 
s 	�      F  , , 
s f 
s . ; . ; f 
s f      F  , , � � � ^ [ ^ [ � � �      F  , ,  &  � � � � &  &      F  , , �  V �  [  [  V �  V      F  , , � f � . [ . [ f � f      F  , , � F �  [  [ F � F      F  , , � 6 � � [ � [ 6 � 6      F  , ,  F   �  � F  F      F  , , �  � � 	� � 	�  �       F  , ,  �  ^ � ^ � �  �      F  , ,  �  � � � � �  �      F  , ,  ��  �� � �� � ��  ��      F  , , � � � � [ � [ � � �      F  , , � v � > [ > [ v � v      F  , , � � � � 	� � 	� � � �      F  , , 
s � 
s ^ ; ^ ; � 
s �      F  , , � � � � [ � [ � � �      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , , �  � � [ � [  �       F  , , � f � . 	� . 	� f � f      F  , , 
s F 
s  ;  ; F 
s F      F  , , � �� � �� [ �� [ �� � ��      F  , ,    � � � �         F  , , � � � � 	� � 	� � � �      F  , , � � � � 	� � 	� � � �      F  , ,  �  N � N � �  �      F  , , 
s � 
s �n ; �n ; � 
s �      F  , , � � � �n [ �n [ � � �      F  , ,  �  �n � �n � �  �      F  , , � � � �n 	� �n 	� � � �      F  , , 
s � 
s �^ ; �^ ; � 
s �      F  , , 
s �� 
s �N ; �N ; �� 
s ��      F  , , � �& � �� [ �� [ �& � �&      F  , , � � � �~ [ �~ [ � � �      F  , , � �v � �> 	� �> 	� �v � �v      F  , , 
s �& 
s �� ; �� ; �& 
s �&      F  , , � �� � �� [ �� [ �� � ��      F  , , � � � �~ 	� �~ 	� � � �      F  , , � �V � � [ � [ �V � �V      F  , ,  �v  �> � �> � �v  �v      F  , , 
s � 
s �~ ; �~ ; � 
s �      F  , , � �� � �N 	� �N 	� �� � ��      F  , , 
s �� 
s �n ; �n ; �� 
s ��      F  , , � �� � �n 	� �n 	� �� � ��      F  , , � �� � �n [ �n [ �� � ��      F  , , � �& � �� 	� �� 	� �& � �&      F  , , � �� � �N [ �N [ �� � ��      F  , , � � � �^ 	� �^ 	� � � �      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , , 
s �V 
s � ; � ; �V 
s �V      F  , , � �� � �� [ �� [ �� � ��      F  , ,  �  �� � �� � �  �      F  , , 
s �� 
s � ; � ; �� 
s ��      F  , ,  �f  �. � �. � �f  �f      F  , , � �F � � [ � [ �F � �F      F  , , � �� � � [ � [ �� � ��      F  , ,  ��  � � � � ��  ��      F  , , � � � �� [ �� [ � � �      F  , ,  �  �� � �� � �  �      F  , ,  ��  �� � �� � ��  ��      F  , , � � � �� [ �� [ � � �      F  , ,  ��  � � � � ��  ��      F  , ,  �  �^ � �^ � �  �      F  , , 
s � 
s �� ; �� ; � 
s �      F  , , � �F � � 	� � 	� �F � �F      F  , , 
s �f 
s �. ; �. ; �f 
s �f      F  , ,  ��  �N � �N � ��  ��      F  , ,  �V  � � � � �V  �V      F  , ,  �6  �� � �� � �6  �6      F  , ,  �&  �� � �� � �&  �&      F  , , � �f � �. 	� �. 	� �f � �f      F  , , 
s �F 
s � ; � ; �F 
s �F      F  , , 
s �v 
s �> ; �> ; �v 
s �v      F  , , � �� � � 	� � 	� �� � ��      F  , , � �� � �� 	� �� 	� �� � ��      F  , , � �� � � 	� � 	� �� � ��      F  , ,  �  �~ � �~ � �  �      F  , , � � � �^ [ �^ [ � � �      F  , , � �f � �. [ �. [ �f � �f      F  , , � �v � �> [ �> [ �v � �v      F  , , 
s �� 
s � ; � ; �� 
s ��      F  , , 
s � 
s �� ; �� ; � 
s �      F  , , � � � �� 	� �� 	� � � �      F  , ,  �F  � � � � �F  �F      F  , , � �V � � 	� � 	� �V � �V      F  , , 
s �6 
s �� ; �� ; �6 
s �6      F  , , � �6 � �� [ �� [ �6 � �6      F  , ,  ��  �� � �� � ��  ��      F  , , � � � �� 	� �� 	� � � �      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , , � �� � �� 	� �� 	� �� � ��      F  , , � �� � � [ � [ �� � ��      F  , , � �6 � �� 	� �� 	� �6 � �6      F  , ,  ��  �n � �n � ��  ��      F  , , 
s Ԗ 
s �^ ; �^ ; Ԗ 
s Ԗ      F  , , � �& � �� 	� �� 	� �& � �&      F  , , � �V � � [ � [ �V � �V      F  , , � ɦ � �n 	� �n 	� ɦ � ɦ      F  , , � ׶ � �~ 	� �~ 	� ׶ � ׶      F  , ,  ��  Ю � Ю � ��  ��      F  , , � �� � Ю [ Ю [ �� � ��      F  , ,  ��  ۞ � ۞ � ��  ��      F  , , � �V � � 	� � 	� �V � �V      F  , , 
s �f 
s �. ; �. ; �f 
s �f      F  , , � ɦ � �n [ �n [ ɦ � ɦ      F  , ,  ɦ  �n � �n � ɦ  ɦ      F  , ,  �&  �� � �� � �&  �&      F  , , � �F � � 	� � 	� �F � �F      F  , , 
s �& 
s �� ; �� ; �& 
s �&      F  , , � �� � ۞ [ ۞ [ �� � ��      F  , ,  ��  ޾ � ޾ � ��  ��      F  , , � �6 � �� 	� �� 	� �6 � �6      F  , ,  �  �� � �� � �  �      F  , , � �f � �. 	� �. 	� �f � �f      F  , ,  ��  ͎ � ͎ � ��  ��      F  , , � ߆ � �N [ �N [ ߆ � ߆      F  , , 
s � 
s �� ; �� ; � 
s �      F  , , � ׶ � �~ [ �~ [ ׶ � ׶      F  , , � �& � �� [ �� [ �& � �&      F  , , 
s �6 
s �� ; �� ; �6 
s �6      F  , , � �� � ޾ [ ޾ [ �� � ��      F  , , � �6 � �� [ �� [ �6 � �6      F  , , � �� � ͎ [ ͎ [ �� � ��      F  , ,  ߆  �N � �N � ߆  ߆      F  , ,  �F  � � � � �F  �F      F  , , � ߆ � �N 	� �N 	� ߆ � ߆      F  , , � �� � Ю 	� Ю 	� �� � ��      F  , ,  Ԗ  �^ � �^ � Ԗ  Ԗ      F  , , � �f � �. [ �. [ �f � �f      F  , , 
s �v 
s �> ; �> ; �v 
s �v      F  , , � � � �� [ �� [ � � �      F  , ,  ׶  �~ � �~ � ׶  ׶      F  , , 
s �� 
s ޾ ; ޾ ; �� 
s ��      F  , ,  �  �� � �� � �  �      F  , ,  �v  �> � �> � �v  �v      F  , , 
s � 
s �� ; �� ; � 
s �      F  , , � �� � ޾ 	� ޾ 	� �� � ��      F  , , � � � �� 	� �� 	� � � �      F  , , � Ԗ � �^ 	� �^ 	� Ԗ � Ԗ      F  , , 
s ׶ 
s �~ ; �~ ; ׶ 
s ׶      F  , , 
s �� 
s ۞ ; ۞ ; �� 
s ��      F  , ,  �f  �. � �. � �f  �f      F  , , � � � �� [ �� [ � � �      F  , ,  �6  �� � �� � �6  �6      F  , ,  �  �� � �� � �  �      F  , , 
s � 
s �� ; �� ; � 
s �      F  , ,  �V  � � � � �V  �V      F  , , � Ԗ � �^ [ �^ [ Ԗ � Ԗ      F  , , � �F � � [ � [ �F � �F      F  , , 
s �V 
s � ; � ; �V 
s �V      F  , , 
s ɦ 
s �n ; �n ; ɦ 
s ɦ      F  , , � � � �� [ �� [ � � �      F  , , 
s �� 
s ͎ ; ͎ ; �� 
s ��      F  , , � �� � ۞ 	� ۞ 	� �� � ��      F  , , 
s �F 
s � ; � ; �F 
s �F      F  , , � �� � ͎ 	� ͎ 	� �� � ��      F  , , 
s �� 
s Ю ; Ю ; �� 
s ��      F  , , � �v � �> 	� �> 	� �v � �v      F  , , � �v � �> [ �> [ �v � �v      F  , , � � � �� 	� �� 	� � � �      F  , , 
s ߆ 
s �N ; �N ; ߆ 
s ߆      F  , , � � � �� 	� �� 	� � � �      F  , ,  �� 3�  �� 4�  �� 4�  �� 3�  �� 3�      F  , ,  �K 3�  �K 4�  � 4�  � 3�  �K 3�      F  , ,  �� 3�  �� 4�  �� 4�  �� 3�  �� 3�      F  , ,  �+ 3�  �+ 4�  �� 4�  �� 3�  �+ 3�      F  , ,  �� �&  �� ��  �� ��  �� �&  �� �&      F  , ,  �� �&  �� ��  �� ��  �� �&  �� �&      F  , ,  �K �&  �K ��  � ��  � �&  �K �&      F  , ,  �+ �&  �+ ��  �� ��  �� �&  �+ �&      F  , ,  �� �f  �� �.  �� �.  �� �f  �� �f      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �� �6  �� ��  �� ��  �� �6  �� �6      F  , ,  �� �F  �� �  �� �  �� �F  �� �F      F  , ,  �� ��  �� �n  �� �n  �� ��  �� ��      F  , ,  �� ��  �� �~  �� �~  �� ��  �� ��      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� ��  �� �N  �� �N  �� ��  �� ��      F  , ,  �� ��  �� �N  �� �N  �� ��  �� ��      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �� �f  �� �.  �� �.  �� �f  �� �f      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �� �F  �� �  �� �  �� �F  �� �F      F  , ,  �� ��  �� �~  �� �~  �� ��  �� ��      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �K ��  �K �~  � �~  � ��  �K ��      F  , ,  �K �&  �K ��  � ��  � �&  �K �&      F  , ,  �K ��  �K �^  � �^  � ��  �K ��      F  , ,  �K �  �K ��  � ��  � �  �K �      F  , ,  �K �v  �K �>  � �>  � �v  �K �v      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �K �V  �K �  � �  � �V  �K �V      F  , ,  �+ ��  �+ �~  �� �~  �� ��  �+ ��      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �+ �&  �+ ��  �� ��  �� �&  �+ �&      F  , ,  �K �6  �K ��  � ��  � �6  �K �6      F  , ,  �+ ��  �+ �^  �� �^  �� ��  �+ ��      F  , ,  �K ��  �K �n  � �n  � ��  �K ��      F  , ,  �+ �  �+ ��  �� ��  �� �  �+ �      F  , ,  �K �  �K ��  � ��  � �  �K �      F  , ,  �+ �v  �+ �>  �� �>  �� �v  �+ �v      F  , ,  �K ��  �K �N  � �N  � ��  �K ��      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �+ �V  �+ �  �� �  �� �V  �+ �V      F  , ,  �� �v  �� �>  �� �>  �� �v  �� �v      F  , ,  �K �f  �K �.  � �.  � �f  �K �f      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �+ �6  �+ ��  �� ��  �� �6  �+ �6      F  , ,  �K �F  �K �  � �  � �F  �K �F      F  , ,  �+ ��  �+ �n  �� �n  �� ��  �+ ��      F  , ,  �K ��  �K �~  � �~  � ��  �K ��      F  , ,  �+ �  �+ ��  �� ��  �� �  �+ �      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �+ ��  �+ �N  �� �N  �� ��  �+ ��      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �+ �f  �+ �.  �� �.  �� �f  �+ �f      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �+ �F  �+ �  �� �  �� �F  �+ �F      F  , ,  �� ��  �� �~  �� �~  �� ��  �� ��      F  , ,  �+ ��  �+ �~  �� �~  �� ��  �+ ��      F  , ,  �� �&  �� ��  �� ��  �� �&  �� �&      F  , ,  �� �V  �� �  �� �  �� �V  �� �V      F  , ,  �� ��  �� �^  �� �^  �� ��  �� ��      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� �v  �� �>  �� �>  �� �v  �� �v      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �� �V  �� �  �� �  �� �V  �� �V      F  , ,  �� ��  �� �~  �� �~  �� ��  �� ��      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �� �&  �� ��  �� ��  �� �&  �� �&      F  , ,  �� �6  �� ��  �� ��  �� �6  �� �6      F  , ,  �� ��  �� �^  �� �^  �� ��  �� ��      F  , ,  �� ��  �� �n  �� �n  �� ��  �� ��      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� oF  �� p  �� p  �� oF  �� oF      F  , ,  �+ p�  �+ q�  �� q�  �� p�  �+ p�      F  , ,  �� {�  �� |�  �� |�  �� {�  �� {�      F  , ,  �� m�  �� n~  �� n~  �� m�  �� m�      F  , ,  �� z6  �� z�  �� z�  �� z6  �� z6      F  , ,  �+ u�  �+ vN  �� vN  �� u�  �+ u�      F  , ,  �� l&  �� l�  �� l�  �� l&  �� l&      F  , ,  �+ w  �+ w�  �� w�  �� w  �+ w      F  , ,  �� x�  �� yn  �� yn  �� x�  �� x�      F  , ,  �� j�  �� k^  �� k^  �� j�  �� j�      F  , ,  �� ��  �� �^  �� �^  �� ��  �� ��      F  , ,  �� w  �� w�  �� w�  �� w  �� w      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� u�  �� vN  �� vN  �� u�  �� u�      F  , ,  �� �v  �� �>  �� �>  �� �v  �� �v      F  , ,  �� s�  �� t�  �� t�  �� s�  �� s�      F  , ,  �� rf  �� s.  �� s.  �� rf  �� rf      F  , ,  �� ~�  �� �  �� �  �� ~�  �� ~�      F  , ,  �� p�  �� q�  �� q�  �� p�  �� p�      F  , ,  �� }V  �� ~  �� ~  �� }V  �� }V      F  , ,  �+ l&  �+ l�  �� l�  �� l&  �+ l&      F  , ,  �� oF  �� p  �� p  �� oF  �� oF      F  , ,  �� {�  �� |�  �� |�  �� {�  �� {�      F  , ,  �K ��  �K �^  � �^  � ��  �K ��      F  , ,  �+ rf  �+ s.  �� s.  �� rf  �+ rf      F  , ,  �K �  �K ��  � ��  � �  �K �      F  , ,  �� m�  �� n~  �� n~  �� m�  �� m�      F  , ,  �K �v  �K �>  � �>  � �v  �K �v      F  , ,  �� z6  �� z�  �� z�  �� z6  �� z6      F  , ,  �K ~�  �K �  � �  � ~�  �K ~�      F  , ,  �� l&  �� l�  �� l�  �� l&  �� l&      F  , ,  �K }V  �K ~  � ~  � }V  �K }V      F  , ,  �� ��  �� �^  �� �^  �� ��  �� ��      F  , ,  �� j�  �� k^  �� k^  �� j�  �� j�      F  , ,  �K {�  �K |�  � |�  � {�  �K {�      F  , ,  �� x�  �� yn  �� yn  �� x�  �� x�      F  , ,  �+ j�  �+ k^  �� k^  �� j�  �+ j�      F  , ,  �K z6  �K z�  � z�  � z6  �K z6      F  , ,  �� w  �� w�  �� w�  �� w  �� w      F  , ,  �K l&  �K l�  � l�  � l&  �K l&      F  , ,  �+ ��  �+ �^  �� �^  �� ��  �+ ��      F  , ,  �K x�  �K yn  � yn  � x�  �K x�      F  , ,  �+ oF  �+ p  �� p  �� oF  �+ oF      F  , ,  �+ �  �+ ��  �� ��  �� �  �+ �      F  , ,  �K w  �K w�  � w�  � w  �K w      F  , ,  �� u�  �� vN  �� vN  �� u�  �� u�      F  , ,  �+ �v  �+ �>  �� �>  �� �v  �+ �v      F  , ,  �K u�  �K vN  � vN  � u�  �K u�      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �+ ~�  �+ �  �� �  �� ~�  �+ ~�      F  , ,  �K s�  �K t�  � t�  � s�  �K s�      F  , ,  �� s�  �� t�  �� t�  �� s�  �� s�      F  , ,  �+ }V  �+ ~  �� ~  �� }V  �+ }V      F  , ,  �+ s�  �+ t�  �� t�  �� s�  �+ s�      F  , ,  �K rf  �K s.  � s.  � rf  �K rf      F  , ,  �� �v  �� �>  �� �>  �� �v  �� �v      F  , ,  �+ {�  �+ |�  �� |�  �� {�  �+ {�      F  , ,  �� rf  �� s.  �� s.  �� rf  �� rf      F  , ,  �K p�  �K q�  � q�  � p�  �K p�      F  , ,  �K j�  �K k^  � k^  � j�  �K j�      F  , ,  �+ z6  �+ z�  �� z�  �� z6  �+ z6      F  , ,  �� ~�  �� �  �� �  �� ~�  �� ~�      F  , ,  �K oF  �K p  � p  � oF  �K oF      F  , ,  �� p�  �� q�  �� q�  �� p�  �� p�      F  , ,  �+ x�  �+ yn  �� yn  �� x�  �+ x�      F  , ,  �+ m�  �+ n~  �� n~  �� m�  �+ m�      F  , ,  �K m�  �K n~  � n~  � m�  �K m�      F  , ,  �� }V  �� ~  �� ~  �� }V  �� }V      F  , ,  �K Nv  �K O>  � O>  � Nv  �K Nv      F  , ,  �� Nv  �� O>  �� O>  �� Nv  �� Nv      F  , ,  �� Nv  �� O>  �� O>  �� Nv  �� Nv      F  , ,  �+ Nv  �+ O>  �� O>  �� Nv  �+ Nv      F  , ,  �K S&  �K S�  � S�  � S&  �K S&      F  , ,  �� \�  �� ]N  �� ]N  �� \�  �� \�      F  , ,  �+ i  �+ i�  �� i�  �� i  �+ i      F  , ,  �� Z�  �� [�  �� [�  �� Z�  �� Z�      F  , ,  �+ ^  �+ ^�  �� ^�  �� ^  �+ ^      F  , ,  �K Q�  �K R^  � R^  � Q�  �K Q�      F  , ,  �� Yf  �� Z.  �� Z.  �� Yf  �� Yf      F  , ,  �K P  �K P�  � P�  � P  �K P      F  , ,  �+ \�  �+ ]N  �� ]N  �� \�  �+ \�      F  , ,  �� W�  �� X�  �� X�  �� W�  �� W�      F  , ,  �K ^  �K ^�  � ^�  � ^  �K ^      F  , ,  �� i  �� i�  �� i�  �� i  �� i      F  , ,  �K T�  �K U~  � U~  � T�  �K T�      F  , ,  �� VF  �� W  �� W  �� VF  �� VF      F  , ,  �+ gv  �+ h>  �� h>  �� gv  �+ gv      F  , ,  �� gv  �� h>  �� h>  �� gv  �� gv      F  , ,  �� T�  �� U~  �� U~  �� T�  �� T�      F  , ,  �+ Z�  �+ [�  �� [�  �� Z�  �+ Z�      F  , ,  �� S&  �� S�  �� S�  �� S&  �� S&      F  , ,  �� e�  �� f�  �� f�  �� e�  �� e�      F  , ,  �� Q�  �� R^  �� R^  �� Q�  �� Q�      F  , ,  �� dV  �� e  �� e  �� dV  �� dV      F  , ,  �K \�  �K ]N  � ]N  � \�  �K \�      F  , ,  �� P  �� P�  �� P�  �� P  �� P      F  , ,  �+ Yf  �+ Z.  �� Z.  �� Yf  �+ Yf      F  , ,  �� b�  �� c�  �� c�  �� b�  �� b�      F  , ,  �K b�  �K c�  � c�  � b�  �K b�      F  , ,  �K _�  �K `n  � `n  � _�  �K _�      F  , ,  �� a6  �� a�  �� a�  �� a6  �� a6      F  , ,  �+ e�  �+ f�  �� f�  �� e�  �+ e�      F  , ,  �� _�  �� `n  �� `n  �� _�  �� _�      F  , ,  �+ W�  �+ X�  �� X�  �� W�  �+ W�      F  , ,  �� ^  �� ^�  �� ^�  �� ^  �� ^      F  , ,  �K e�  �K f�  � f�  � e�  �K e�      F  , ,  �K Z�  �K [�  � [�  � Z�  �K Z�      F  , ,  �� \�  �� ]N  �� ]N  �� \�  �� \�      F  , ,  �K i  �K i�  � i�  � i  �K i      F  , ,  �� Z�  �� [�  �� [�  �� Z�  �� Z�      F  , ,  �+ VF  �+ W  �� W  �� VF  �+ VF      F  , ,  �+ dV  �+ e  �� e  �� dV  �+ dV      F  , ,  �� Yf  �� Z.  �� Z.  �� Yf  �� Yf      F  , ,  �K Yf  �K Z.  � Z.  � Yf  �K Yf      F  , ,  �� i  �� i�  �� i�  �� i  �� i      F  , ,  �� W�  �� X�  �� X�  �� W�  �� W�      F  , ,  �+ T�  �+ U~  �� U~  �� T�  �+ T�      F  , ,  �K gv  �K h>  � h>  � gv  �K gv      F  , ,  �� VF  �� W  �� W  �� VF  �� VF      F  , ,  �� gv  �� h>  �� h>  �� gv  �� gv      F  , ,  �+ S&  �+ S�  �� S�  �� S&  �+ S&      F  , ,  �� T�  �� U~  �� U~  �� T�  �� T�      F  , ,  �K W�  �K X�  � X�  � W�  �K W�      F  , ,  �� e�  �� f�  �� f�  �� e�  �� e�      F  , ,  �� S&  �� S�  �� S�  �� S&  �� S&      F  , ,  �+ Q�  �+ R^  �� R^  �� Q�  �+ Q�      F  , ,  �+ b�  �+ c�  �� c�  �� b�  �+ b�      F  , ,  �� Q�  �� R^  �� R^  �� Q�  �� Q�      F  , ,  �� dV  �� e  �� e  �� dV  �� dV      F  , ,  �K a6  �K a�  � a�  � a6  �K a6      F  , ,  �� P  �� P�  �� P�  �� P  �� P      F  , ,  �+ P  �+ P�  �� P�  �� P  �+ P      F  , ,  �� b�  �� c�  �� c�  �� b�  �� b�      F  , ,  �+ _�  �+ `n  �� `n  �� _�  �+ _�      F  , ,  �K VF  �K W  � W  � VF  �K VF      F  , ,  �� a6  �� a�  �� a�  �� a6  �� a6      F  , ,  �� ^  �� ^�  �� ^�  �� ^  �� ^      F  , ,  �+ a6  �+ a�  �� a�  �� a6  �+ a6      F  , ,  �K dV  �K e  � e  � dV  �K dV      F  , ,  �� _�  �� `n  �� `n  �� _�  �� _�      F  , ,  �+ I�  �+ J�  �� J�  �� I�  �+ I�      F  , ,  �+ KV  �+ L  �� L  �� KV  �+ KV      F  , ,  �� H6  �� H�  �� H�  �� H6  �� H6      F  , ,  �+ :&  �+ :�  �� :�  �� :&  �+ :&      F  , ,  �+ E  �+ E�  �� E�  �� E  �+ E      F  , ,  �K :&  �K :�  � :�  � :&  �K :&      F  , ,  �� :&  �� :�  �� :�  �� :&  �� :&      F  , ,  �� F�  �� Gn  �� Gn  �� F�  �� F�      F  , ,  �+ 8�  �+ 9^  �� 9^  �� 8�  �+ 8�      F  , ,  �K H6  �K H�  � H�  � H6  �K H6      F  , ,  �� ;�  �� <~  �� <~  �� ;�  �� ;�      F  , ,  �� E  �� E�  �� E�  �� E  �� E      F  , ,  �K 7  �K 7�  � 7�  � 7  �K 7      F  , ,  �� 7  �� 7�  �� 7�  �� 7  �� 7      F  , ,  �+ 7  �+ 7�  �� 7�  �� 7  �+ 7      F  , ,  �� C�  �� DN  �� DN  �� C�  �� C�      F  , ,  �+ C�  �+ DN  �� DN  �� C�  �+ C�      F  , ,  �� 7  �� 7�  �� 7�  �� 7  �� 7      F  , ,  �� :&  �� :�  �� :�  �� :&  �� :&      F  , ,  �K F�  �K Gn  � Gn  � F�  �K F�      F  , ,  �� A�  �� B�  �� B�  �� A�  �� A�      F  , ,  �+ 5v  �+ 6>  �� 6>  �� 5v  �+ 5v      F  , ,  �� H6  �� H�  �� H�  �� H6  �� H6      F  , ,  �� E  �� E�  �� E�  �� E  �� E      F  , ,  �+ H6  �+ H�  �� H�  �� H6  �+ H6      F  , ,  �� >�  �� ?�  �� ?�  �� >�  �� >�      F  , ,  �� @f  �� A.  �� A.  �� @f  �� @f      F  , ,  �+ A�  �+ B�  �� B�  �� A�  �+ A�      F  , ,  �K E  �K E�  � E�  � E  �K E      F  , ,  �K L�  �K M�  � M�  � L�  �K L�      F  , ,  �� C�  �� DN  �� DN  �� C�  �� C�      F  , ,  �� ;�  �� <~  �� <~  �� ;�  �� ;�      F  , ,  �� 5v  �� 6>  �� 6>  �� 5v  �� 5v      F  , ,  �+ L�  �+ M�  �� M�  �� L�  �+ L�      F  , ,  �K C�  �K DN  � DN  � C�  �K C�      F  , ,  �+ @f  �+ A.  �� A.  �� @f  �+ @f      F  , ,  �K 5v  �K 6>  � 6>  � 5v  �K 5v      F  , ,  �� 5v  �� 6>  �� 6>  �� 5v  �� 5v      F  , ,  �K ;�  �K <~  � <~  � ;�  �K ;�      F  , ,  �K A�  �K B�  � B�  � A�  �K A�      F  , ,  �+ F�  �+ Gn  �� Gn  �� F�  �+ F�      F  , ,  �+ >�  �+ ?�  �� ?�  �� >�  �+ >�      F  , ,  �K KV  �K L  � L  � KV  �K KV      F  , ,  �K 8�  �K 9^  � 9^  � 8�  �K 8�      F  , ,  �K @f  �K A.  � A.  � @f  �K @f      F  , ,  �� L�  �� M�  �� M�  �� L�  �� L�      F  , ,  �� 8�  �� 9^  �� 9^  �� 8�  �� 8�      F  , ,  �+ =F  �+ >  �� >  �� =F  �+ =F      F  , ,  �� A�  �� B�  �� B�  �� A�  �� A�      F  , ,  �� F�  �� Gn  �� Gn  �� F�  �� F�      F  , ,  �� KV  �� L  �� L  �� KV  �� KV      F  , ,  �� 8�  �� 9^  �� 9^  �� 8�  �� 8�      F  , ,  �K >�  �K ?�  � ?�  � >�  �K >�      F  , ,  �� >�  �� ?�  �� ?�  �� >�  �� >�      F  , ,  �� I�  �� J�  �� J�  �� I�  �� I�      F  , ,  �� L�  �� M�  �� M�  �� L�  �� L�      F  , ,  �� @f  �� A.  �� A.  �� @f  �� @f      F  , ,  �� =F  �� >  �� >  �� =F  �� =F      F  , ,  �� I�  �� J�  �� J�  �� I�  �� I�      F  , ,  �+ ;�  �+ <~  �� <~  �� ;�  �+ ;�      F  , ,  �� KV  �� L  �� L  �� KV  �� KV      F  , ,  �K =F  �K >  � >  � =F  �K =F      F  , ,  �� =F  �� >  �� >  �� =F  �� =F      F  , ,  �K I�  �K J�  � J�  � I�  �K I�      F  , ,  �+ �6  �+ ��  �� ��  �� �6  �+ �6      F  , ,  �� �6  �� ��  �� ��  �� �6  �� �6      F  , ,  �� �6  �� ��  �� ��  �� �6  �� �6      F  , ,  �K �6  �K ��  � ��  � �6  �K �6      F  , ,  �+   �+ �  �� �  ��   �+       F  , ,  �� *�  �� +N  �� +N  �� *�  �� *�      F  , ,  �� (�  �� )�  �� )�  �� (�  �� (�      F  , ,  �� 'f  �� (.  �� (.  �� 'f  �� 'f      F  , ,  �+ $F  �+ %  �� %  �� $F  �+ $F      F  , ,  �K 2V  �K 3  � 3  � 2V  �K 2V      F  , ,  �� 2V  �� 3  �� 3  �� 2V  �� 2V      F  , ,  �K 0�  �K 1�  � 1�  � 0�  �K 0�      F  , ,  �� 0�  �� 1�  �� 1�  �� 0�  �� 0�      F  , ,  �� %�  �� &�  �� &�  �� %�  �� %�      F  , ,  �+ v  �+ >  �� >  �� v  �+ v      F  , ,  �+ !&  �+ !�  �� !�  �� !&  �+ !&      F  , ,  �K /6  �K /�  � /�  � /6  �K /6      F  , ,  �� /6  �� /�  �� /�  �� /6  �� /6      F  , ,  �� $F  �� %  �� %  �� $F  �� $F      F  , ,  �K -�  �K .n  � .n  � -�  �K -�      F  , ,  �� -�  �� .n  �� .n  �� -�  �� -�      F  , ,  �+ %�  �+ &�  �� &�  �� %�  �+ %�      F  , ,  �K ,  �K ,�  � ,�  � ,  �K ,      F  , ,  �� ,  �� ,�  �� ,�  �� ,  �� ,      F  , ,  �� "�  �� #~  �� #~  �� "�  �� "�      F  , ,  �K *�  �K +N  � +N  � *�  �K *�      F  , ,  �� *�  �� +N  �� +N  �� *�  �� *�      F  , ,  �K (�  �K )�  � )�  � (�  �K (�      F  , ,  �� (�  �� )�  �� )�  �� (�  �� (�      F  , ,  �+ �  �+ �  �� �  �� �  �+ �      F  , ,  �� !&  �� !�  �� !�  �� !&  �� !&      F  , ,  �K 'f  �K (.  � (.  � 'f  �K 'f      F  , ,  �� 'f  �� (.  �� (.  �� 'f  �� 'f      F  , ,  �� �  ��  ^  ��  ^  �� �  �� �      F  , ,  �K %�  �K &�  � &�  � %�  �K %�      F  , ,  �� %�  �� &�  �� &�  �� %�  �� %�      F  , ,  �K $F  �K %  � %  � $F  �K $F      F  , ,  �� $F  �� %  �� %  �� $F  �� $F      F  , ,  �K "�  �K #~  � #~  � "�  �K "�      F  , ,  �� "�  �� #~  �� #~  �� "�  �� "�      F  , ,  ��   �� �  �� �  ��   ��       F  , ,  �� 2V  �� 3  �� 3  �� 2V  �� 2V      F  , ,  �K !&  �K !�  � !�  � !&  �K !&      F  , ,  �� !&  �� !�  �� !�  �� !&  �� !&      F  , ,  �+ �  �+  ^  ��  ^  �� �  �+ �      F  , ,  �� ,  �� ,�  �� ,�  �� ,  �� ,      F  , ,  �K �  �K  ^  �  ^  � �  �K �      F  , ,  �� �  ��  ^  ��  ^  �� �  �� �      F  , ,  �� v  �� >  �� >  �� v  �� v      F  , ,  �K v  �K >  � >  � v  �K v      F  , ,  �� 0�  �� 1�  �� 1�  �� 0�  �� 0�      F  , ,  �K   �K �  � �  �   �K       F  , ,  ��   �� �  �� �  ��   ��       F  , ,  �+ V  �+   ��   �� V  �+ V      F  , ,  �� v  �� >  �� >  �� v  �� v      F  , ,  �+ 2V  �+ 3  �� 3  �� 2V  �+ 2V      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �K �  �K �  � �  � �  �K �      F  , ,  �� V  ��   ��   �� V  �� V      F  , ,  �+ 0�  �+ 1�  �� 1�  �� 0�  �+ 0�      F  , ,  �� /6  �� /�  �� /�  �� /6  �� /6      F  , ,  �+ /6  �+ /�  �� /�  �� /6  �+ /6      F  , ,  �� V  ��   ��   �� V  �� V      F  , ,  �+ -�  �+ .n  �� .n  �� -�  �+ -�      F  , ,  �K V  �K   �   � V  �K V      F  , ,  �+ "�  �+ #~  �� #~  �� "�  �+ "�      F  , ,  �+ 'f  �+ (.  �� (.  �� 'f  �+ 'f      F  , ,  �+ ,  �+ ,�  �� ,�  �� ,  �+ ,      F  , ,  �� -�  �� .n  �� .n  �� -�  �� -�      F  , ,  �+ *�  �+ +N  �� +N  �� *�  �+ *�      F  , ,  �+ (�  �+ )�  �� )�  �� (�  �+ (�      F  , ,  �+ v  �+ >  �� >  �� v  �+ v      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �+ 	�  �+ 
~  �� 
~  �� 	�  �+ 	�      F  , ,  �� v  �� >  �� >  �� v  �� v      F  , ,  �K v  �K >  � >  � v  �K v      F  , ,  �+ �  �+ ^  �� ^  �� �  �+ �      F  , ,  �+ &  �+ �  �� �  �� &  �+ &      F  , ,  �� 	�  �� 
~  �� 
~  �� 	�  �� 	�      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �K �  �K �  � �  � �  �K �      F  , ,  �� 6  �� �  �� �  �� 6  �� 6      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �K �  �K �  � �  � �  �K �      F  , ,  �+ �  �+ �  �� �  �� �  �+ �      F  , ,  ��  V  ��   ��   ��  V  ��  V      F  , ,  �K  V  �K   �   �  V  �K  V      F  , ,  �� �  �� N  �� N  �� �  �� �      F  , ,  �K �  �K N  � N  � �  �K �      F  , ,  �+ �  �+ �  �� �  �� �  �+ �      F  , ,  �� F  ��   ��   �� F  �� F      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �K F  �K   �   � F  �K F      F  , ,  �� �  �� ^  �� ^  �� �  �� �      F  , ,  �+   �+ �  �� �  ��   �+       F  , ,  �K 6  �K �  � �  � 6  �K 6      F  , ,  �� �  �� n  �� n  �� �  �� �      F  , ,  �+ f  �+ .  �� .  �� f  �+ f      F  , ,  �+   �+ �  �� �  ��   �+       F  , ,  �� 	�  �� 
~  �� 
~  �� 	�  �� 	�      F  , ,  �K 	�  �K 
~  � 
~  � 	�  �K 	�      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �K �  �K �  � �  � �  �K �      F  , ,  �K �  �K n  � n  � �  �K �      F  , ,  �+  V  �+   ��   ��  V  �+  V      F  , ,  �� F  ��   ��   �� F  �� F      F  , ,  �� &  �� �  �� �  �� &  �� &      F  , ,  �K &  �K �  � �  � &  �K &      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �+ 6  �+ �  �� �  �� 6  �+ 6      F  , ,  �+ �  �+ n  �� n  �� �  �+ �      F  , ,  �� v  �� >  �� >  �� v  �� v      F  , ,  �+ �  �+ �  �� �  �� �  �+ �      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  ��   �� �  �� �  ��   ��       F  , ,  �� �  �� ^  �� ^  �� �  �� �      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �K �  �K ^  � ^  � �  �K �      F  , ,  �� 6  �� �  �� �  �� 6  �� 6      F  , ,  ��  V  ��   ��   ��  V  ��  V      F  , ,  �� f  �� .  �� .  �� f  �� f      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �� &  �� �  �� �  �� &  �� &      F  , ,  �� �  �� n  �� n  �� �  �� �      F  , ,  �K f  �K .  � .  � f  �K f      F  , ,  ��   �� �  �� �  ��   ��       F  , ,  �+ �  �+ N  �� N  �� �  �+ �      F  , ,  ��   �� �  �� �  ��   ��       F  , ,  �+ F  �+   ��   �� F  �+ F      F  , ,  ��   �� �  �� �  ��   ��       F  , ,  �� �  �� N  �� N  �� �  �� �      F  , ,  �K   �K �  � �  �   �K       F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �K �  �K �  � �  � �  �K �      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �K   �K �  � �  �   �K       F  , ,  �+ �  �+ �  �� �  �� �  �+ �      F  , ,  �� f  �� .  �� .  �� f  �� f      F  , ,  �K �  �K �n  � �n  � �  �K �      F  , ,  �� �  �� �n  �� �n  �� �  �� �      F  , ,  �+ �  �+ �n  �� �n  �� �  �+ �      F  , ,  �� �  �� �n  �� �n  �� �  �� �      F  , ,  �+ �&  �+ ��  �� ��  �� �&  �+ �&      F  , ,  �� �F  �� �  �� �  �� �F  �� �F      F  , ,  �K �v  �K �>  � �>  � �v  �K �v      F  , ,  �� �&  �� ��  �� ��  �� �&  �� �&      F  , ,  �� �f  �� �.  �� �.  �� �f  �� �f      F  , ,  �� �6  �� ��  �� ��  �� �6  �� �6      F  , ,  �+ ��  �+ �  �� �  �� ��  �+ ��      F  , ,  �K ��  �K �  � �  � ��  �K ��      F  , ,  �� ��  �� �  �� �  �� ��  �� ��      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �+ ��  �+ �n  �� �n  �� ��  �+ ��      F  , ,  �� �V  �� �  �� �  �� �V  �� �V      F  , ,  �� �  �� �~  �� �~  �� �  �� �      F  , ,  �+ �V  �+ �  �� �  �� �V  �+ �V      F  , ,  �+ �  �+ ��  �� ��  �� �  �+ �      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� �V  �� �  �� �  �� �V  �� �V      F  , ,  �+ �v  �+ �>  �� �>  �� �v  �+ �v      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �+ �  �+ �^  �� �^  �� �  �+ �      F  , ,  �� �  �� �^  �� �^  �� �  �� �      F  , ,  �� ��  �� �n  �� �n  �� ��  �� ��      F  , ,  �K ��  �K �n  � �n  � ��  �K ��      F  , ,  �K �6  �K ��  � ��  � �6  �K �6      F  , ,  �K �  �K ��  � ��  � �  �K �      F  , ,  �+ ��  �+ �N  �� �N  �� ��  �+ ��      F  , ,  �� ��  �� �N  �� �N  �� ��  �� ��      F  , ,  �+ ��  �+ �  �� �  �� ��  �+ ��      F  , ,  �� ��  �� �n  �� �n  �� ��  �� ��      F  , ,  �� �&  �� ��  �� ��  �� �&  �� �&      F  , ,  �K ��  �K �N  � �N  � ��  �K ��      F  , ,  �� ��  �� �  �� �  �� ��  �� ��      F  , ,  �� ��  �� �N  �� �N  �� ��  �� ��      F  , ,  �+ �  �+ �~  �� �~  �� �  �+ �      F  , ,  �� ��  �� �  �� �  �� ��  �� ��      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �� �  �� �~  �� �~  �� �  �� �      F  , ,  �K �f  �K �.  � �.  � �f  �K �f      F  , ,  �� ��  �� �  �� �  �� ��  �� ��      F  , ,  �+ �6  �+ ��  �� ��  �� �6  �+ �6      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �� �6  �� ��  �� ��  �� �6  �� �6      F  , ,  �K �F  �K �  � �  � �F  �K �F      F  , ,  �+ �  �+ ��  �� ��  �� �  �+ �      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� �v  �� �>  �� �>  �� �v  �� �v      F  , ,  �� �  �� �^  �� �^  �� �  �� �      F  , ,  �K �  �K �~  � �~  � �  �K �      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �� �v  �� �>  �� �>  �� �v  �� �v      F  , ,  �� �F  �� �  �� �  �� �F  �� �F      F  , ,  �+ �f  �+ �.  �� �.  �� �f  �+ �f      F  , ,  �K �&  �K ��  � ��  � �&  �K �&      F  , ,  �K �V  �K �  � �  � �V  �K �V      F  , ,  �� �f  �� �.  �� �.  �� �f  �� �f      F  , ,  �+ �F  �+ �  �� �  �� �F  �+ �F      F  , ,  �K �  �K �^  � �^  � �  �K �      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �K �  �K ��  � ��  � �  �K �      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �K ��  �K �  � �  � ��  �K ��      F  , ,  �K �  �K ��  � ��  � �  �K �      F  , ,  �K ��  �K ޾  � ޾  � ��  �K ��      F  , ,  �� �&  �� ��  �� ��  �� �&  �� �&      F  , ,  �K �&  �K ��  � ��  � �&  �K �&      F  , ,  �� ɦ  �� �n  �� �n  �� ɦ  �� ɦ      F  , ,  �+ �V  �+ �  �� �  �� �V  �+ �V      F  , ,  �� ��  �� Ю  �� Ю  �� ��  �� ��      F  , ,  �+ ׶  �+ �~  �� �~  �� ׶  �+ ׶      F  , ,  �� �V  �� �  �� �  �� �V  �� �V      F  , ,  �� Ԗ  �� �^  �� �^  �� Ԗ  �� Ԗ      F  , ,  �� ߆  �� �N  �� �N  �� ߆  �� ߆      F  , ,  �� �v  �� �>  �� �>  �� �v  �� �v      F  , ,  �+ ��  �+ ͎  �� ͎  �� ��  �+ ��      F  , ,  �+ ��  �+ ۞  �� ۞  �� ��  �+ ��      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� �F  �� �  �� �  �� �F  �� �F      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �K �6  �K ��  � ��  � �6  �K �6      F  , ,  �� ��  �� ۞  �� ۞  �� ��  �� ��      F  , ,  �+ Ԗ  �+ �^  �� �^  �� Ԗ  �+ Ԗ      F  , ,  �+ ��  �+ ޾  �� ޾  �� ��  �+ ��      F  , ,  �� ��  �� ޾  �� ޾  �� ��  �� ��      F  , ,  �� �v  �� �>  �� �>  �� �v  �� �v      F  , ,  �K Ԗ  �K �^  � �^  � Ԗ  �K Ԗ      F  , ,  �K ߆  �K �N  � �N  � ߆  �K ߆      F  , ,  �� ��  �� ޾  �� ޾  �� ��  �� ��      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �+ �6  �+ ��  �� ��  �� �6  �+ �6      F  , ,  �+ ɦ  �+ �n  �� �n  �� ɦ  �+ ɦ      F  , ,  �� ��  �� Ю  �� Ю  �� ��  �� ��      F  , ,  �K �  �K ��  � ��  � �  �K �      F  , ,  �K �v  �K �>  � �>  � �v  �K �v      F  , ,  �� �6  �� ��  �� ��  �� �6  �� �6      F  , ,  �+ �F  �+ �  �� �  �� �F  �+ �F      F  , ,  �� �F  �� �  �� �  �� �F  �� �F      F  , ,  �K �F  �K �  � �  � �F  �K �F      F  , ,  �+ ��  �+ Ю  �� Ю  �� ��  �+ ��      F  , ,  �+ �v  �+ �>  �� �>  �� �v  �+ �v      F  , ,  �� �V  �� �  �� �  �� �V  �� �V      F  , ,  �K �f  �K �.  � �.  � �f  �K �f      F  , ,  �K �  �K ��  � ��  � �  �K �      F  , ,  �+ ߆  �+ �N  �� �N  �� ߆  �+ ߆      F  , ,  �� ׶  �� �~  �� �~  �� ׶  �� ׶      F  , ,  �� ��  �� ۞  �� ۞  �� ��  �� ��      F  , ,  �K ��  �K ۞  � ۞  � ��  �K ��      F  , ,  �+ �  �+ ��  �� ��  �� �  �+ �      F  , ,  �� ��  �� ͎  �� ͎  �� ��  �� ��      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� ��  �� ͎  �� ͎  �� ��  �� ��      F  , ,  �K ��  �K ͎  � ͎  � ��  �K ��      F  , ,  �+ �&  �+ ��  �� ��  �� �&  �+ �&      F  , ,  �� ׶  �� �~  �� �~  �� ׶  �� ׶      F  , ,  �� �6  �� ��  �� ��  �� �6  �� �6      F  , ,  �+ �  �+ ��  �� ��  �� �  �+ �      F  , ,  �K ɦ  �K �n  � �n  � ɦ  �K ɦ      F  , ,  �� Ԗ  �� �^  �� �^  �� Ԗ  �� Ԗ      F  , ,  �K ׶  �K �~  � �~  � ׶  �K ׶      F  , ,  �� ߆  �� �N  �� �N  �� ߆  �� ߆      F  , ,  �K ��  �K Ю  � Ю  � ��  �K ��      F  , ,  �� ɦ  �� �n  �� �n  �� ɦ  �� ɦ      F  , ,  �� �f  �� �.  �� �.  �� �f  �� �f      F  , ,  �� �&  �� ��  �� ��  �� �&  �� �&      F  , ,  �K �V  �K �  � �  � �V  �K �V      F  , ,  �+ �f  �+ �.  �� �.  �� �f  �+ �f      F  , ,  �+ �  �+ ��  �� ��  �� �  �+ �      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� �f  �� �.  �� �.  �� �f  �� �f      F  , ,  �+ Z�  �+ [~  �� [~  �� Z�  �+ Z�      F  , ,  �K Z�  �K [~  � [~  � Z�  �K Z�      F  , ,  �� Z�  �� [~  �� [~  �� Z�  �� Z�      F  , ,  �� Z�  �� [~  �� [~  �� Z�  �� Z�      F  , ,  �� �f  �� �.  �� �.  �� �f  �� �f      F  , ,  �+ �f  �+ �.  �� �.  �� �f  �+ �f      F  , ,  �K �f  �K �.  � �.  � �f  �K �f      F  , ,  �� �f  �� �.  �� �.  �� �f  �� �f      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �K �6  �K ��  � ��  � �6  �K �6      F  , ,  �� �f  �� �.  �� �.  �� �f  �� �f      F  , ,  �K �V  �K �  � �  � �V  �K �V      F  , ,  �K ��  �K �n  � �n  � ��  �K ��      F  , ,  �� ��  �� �^  �� �^  �� ��  �� ��      F  , ,  �K �  �K ��  � ��  � �  �K �      F  , ,  �K ��  �K �N  � �N  � ��  �K ��      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� ��  ��   ��   �� ��  �� ��      F  , ,  �+ Ɔ  �+ �N  �� �N  �� Ɔ  �+ Ɔ      F  , ,  �� �v  �� �>  �� �>  �� �v  �� �v      F  , ,  �+ ��  �+ ž  �� ž  �� ��  �+ ��      F  , ,  �K Ɔ  �K �N  � �N  � Ɔ  �K Ɔ      F  , ,  �+ �f  �+ �.  �� �.  �� �f  �+ �f      F  , ,  �K ��  �K ž  � ž  � ��  �K ��      F  , ,  �� Ɔ  �� �N  �� �N  �� Ɔ  �� Ɔ      F  , ,  �+ ��  �+   ��   �� ��  �+ ��      F  , ,  �� ��  �� ž  �� ž  �� ��  �� ��      F  , ,  �+ �F  �+ �  �� �  �� �F  �+ �F      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �K �f  �K �.  � �.  � �f  �K �f      F  , ,  �� �f  �� �.  �� �.  �� �f  �� �f      F  , ,  �+ ��  �+ �~  �� �~  �� ��  �+ ��      F  , ,  �K ��  �K   �   � ��  �K ��      F  , ,  �� ��  ��   ��   �� ��  �� ��      F  , ,  �+ �&  �+ ��  �� ��  �� �&  �+ �&      F  , ,  �� �F  �� �  �� �  �� �F  �� �F      F  , ,  �+ ��  �+ �^  �� �^  �� ��  �+ ��      F  , ,  �� �V  �� �  �� �  �� �V  �� �V      F  , ,  �K �F  �K �  � �  � �F  �K �F      F  , ,  �� ��  �� �~  �� �~  �� ��  �� ��      F  , ,  �� �F  �� �  �� �  �� �F  �� �F      F  , ,  �+ �  �+ ��  �� ��  �� �  �+ �      F  , ,  �K ��  �K �~  � �~  � ��  �K ��      F  , ,  �� �&  �� ��  �� ��  �� �&  �� �&      F  , ,  �+ �v  �+ �>  �� �>  �� �v  �+ �v      F  , ,  �� ��  �� �^  �� �^  �� ��  �� ��      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �� ��  �� ž  �� ž  �� ��  �� ��      F  , ,  �K �&  �K ��  � ��  � �&  �K �&      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �+ �V  �+ �  �� �  �� �V  �+ �V      F  , ,  �� �v  �� �>  �� �>  �� �v  �� �v      F  , ,  �K ��  �K �^  � �^  � ��  �K ��      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �+ �6  �+ ��  �� ��  �� �6  �+ �6      F  , ,  �� �V  �� �  �� �  �� �V  �� �V      F  , ,  �+ ��  �+ �n  �� �n  �� ��  �+ ��      F  , ,  �K �  �K ��  � ��  � �  �K �      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �+ �  �+ ��  �� ��  �� �  �+ �      F  , ,  �� �6  �� ��  �� ��  �� �6  �� �6      F  , ,  �� �6  �� ��  �� ��  �� �6  �� �6      F  , ,  �+ ��  �+ �N  �� �N  �� ��  �+ ��      F  , ,  �� ��  �� �~  �� �~  �� ��  �� ��      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� ��  �� �n  �� �n  �� ��  �� ��      F  , ,  �K �v  �K �>  � �>  � �v  �K �v      F  , ,  �� Ɔ  �� �N  �� �N  �� Ɔ  �� Ɔ      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� ��  �� �n  �� �n  �� ��  �� ��      F  , ,  �� ��  �� �N  �� �N  �� ��  �� ��      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �� ��  �� �N  �� �N  �� ��  �� ��      F  , ,  �� �&  �� ��  �� ��  �� �&  �� �&      F  , ,  �K ��  �K �~  � �~  � ��  �K ��      F  , ,  �� �F  �� �  �� �  �� �F  �� �F      F  , ,  �� �&  �� ��  �� ��  �� �&  �� �&      F  , ,  �� �V  �� �  �� �  �� �V  �� �V      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �� ��  �� �^  �� �^  �� ��  �� ��      F  , ,  �� �6  �� ��  �� ��  �� �6  �� �6      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �K �&  �K ��  � ��  � �&  �K �&      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �K �6  �K ��  � ��  � �6  �K �6      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �� �F  �� �  �� �  �� �F  �� �F      F  , ,  �+ ��  �+ �^  �� �^  �� ��  �+ ��      F  , ,  �+ ��  �+ �N  �� �N  �� ��  �+ ��      F  , ,  �K ��  �K �n  � �n  � ��  �K ��      F  , ,  �K �f  �K �.  � �.  � �f  �K �f      F  , ,  �K ��  �K �^  � �^  � ��  �K ��      F  , ,  �+ �&  �+ ��  �� ��  �� �&  �+ �&      F  , ,  �� �6  �� ��  �� ��  �� �6  �� �6      F  , ,  �K �  �K ��  � ��  � �  �K �      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �+ �v  �+ �>  �� �>  �� �v  �+ �v      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �K ��  �K �N  � �N  � ��  �K ��      F  , ,  �� ��  �� �~  �� �~  �� ��  �� ��      F  , ,  �� ��  �� �N  �� �N  �� ��  �� ��      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �� ��  �� �n  �� �n  �� ��  �� ��      F  , ,  �K �  �K ��  � ��  � �  �K �      F  , ,  �� ��  �� �^  �� �^  �� ��  �� ��      F  , ,  �+ �6  �+ ��  �� ��  �� �6  �+ �6      F  , ,  �+ �  �+ ��  �� ��  �� �  �+ �      F  , ,  �+ �  �+ ��  �� ��  �� �  �+ �      F  , ,  �� �v  �� �>  �� �>  �� �v  �� �v      F  , ,  �K �v  �K �>  � �>  � �v  �K �v      F  , ,  �+ �V  �+ �  �� �  �� �V  �+ �V      F  , ,  �� �V  �� �  �� �  �� �V  �� �V      F  , ,  �K �F  �K �  � �  � �F  �K �F      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� ��  �� �n  �� �n  �� ��  �� ��      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �+ �f  �+ �.  �� �.  �� �f  �+ �f      F  , ,  �� �&  �� ��  �� ��  �� �&  �� �&      F  , ,  �+ ��  �+ �n  �� �n  �� ��  �+ ��      F  , ,  �� ��  �� �N  �� �N  �� ��  �� ��      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �� �f  �� �.  �� �.  �� �f  �� �f      F  , ,  �+ ��  �+ �~  �� �~  �� ��  �+ ��      F  , ,  �+ �F  �+ �  �� �  �� �F  �+ �F      F  , ,  �� ��  �� �~  �� �~  �� ��  �� ��      F  , ,  �K �V  �K �  � �  � �V  �K �V      F  , ,  �� �v  �� �>  �� �>  �� �v  �� �v      F  , ,  �� �f  �� �.  �� �.  �� �f  �� �f      F  , ,  �� }  �� }�  �� }�  �� }  �� }      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �� �6  �� ��  �� ��  �� �6  �� �6      F  , ,  �� {�  �� |N  �� |N  �� {�  �� {�      F  , ,  �K xf  �K y.  � y.  � xf  �K xf      F  , ,  �+ {�  �+ |N  �� |N  �� {�  �+ {�      F  , ,  �� �  �� ��  �� ��  �� �  �� �      F  , ,  �+ �V  �+ �  �� �  �� �V  �+ �V      F  , ,  �� �F  �� �  �� �  �� �F  �� �F      F  , ,  �� y�  �� z�  �� z�  �� y�  �� y�      F  , ,  �� �v  �� �>  �� �>  �� �v  �� �v      F  , ,  �� ~�  �� n  �� n  �� ~�  �� ~�      F  , ,  �+ y�  �+ z�  �� z�  �� y�  �+ y�      F  , ,  �� xf  �� y.  �� y.  �� xf  �� xf      F  , ,  �� ��  �� �~  �� �~  �� ��  �� ��      F  , ,  �K {�  �K |N  � |N  � {�  �K {�      F  , ,  �� �v  �� �>  �� �>  �� �v  �� �v      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �� }  �� }�  �� }�  �� }  �� }      F  , ,  �� v�  �� w�  �� w�  �� v�  �� v�      F  , ,  �+ xf  �+ y.  �� y.  �� xf  �+ xf      F  , ,  �+ �  �+ ��  �� ��  �� �  �+ �      F  , ,  �� ��  �� �~  �� �~  �� ��  �� ��      F  , ,  �K ~�  �K n  � n  � ~�  �K ~�      F  , ,  �� �V  �� �  �� �  �� �V  �� �V      F  , ,  �� {�  �� |N  �� |N  �� {�  �� {�      F  , ,  �+ v�  �+ w�  �� w�  �� v�  �+ v�      F  , ,  �K �v  �K �>  � �>  � �v  �K �v      F  , ,  �K v�  �K w�  � w�  � v�  �K v�      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �+ �6  �+ ��  �� ��  �� �6  �+ �6      F  , ,  �� y�  �� z�  �� z�  �� y�  �� y�      F  , ,  �K y�  �K z�  � z�  � y�  �K y�      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �K �6  �K ��  � ��  � �6  �K �6      F  , ,  �+ ��  �+ ��  �� ��  �� ��  �+ ��      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �� �&  �� ��  �� ��  �� �&  �� �&      F  , ,  �� �&  �� ��  �� ��  �� �&  �� �&      F  , ,  �K �V  �K �  � �  � �V  �K �V      F  , ,  �+ �v  �+ �>  �� �>  �� �v  �+ �v      F  , ,  �� xf  �� y.  �� y.  �� xf  �� xf      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �� �V  �� �  �� �  �� �V  �� �V      F  , ,  �K ��  �K ��  � ��  � ��  �K ��      F  , ,  �� �F  �� �  �� �  �� �F  �� �F      F  , ,  �+ ~�  �+ n  �� n  �� ~�  �+ ~�      F  , ,  �K �F  �K �  � �  � �F  �K �F      F  , ,  �� �6  �� ��  �� ��  �� �6  �� �6      F  , ,  �+ �&  �+ ��  �� ��  �� �&  �+ �&      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �K ��  �K �~  � �~  � ��  �K ��      F  , ,  �+ �F  �+ �  �� �  �� �F  �+ �F      F  , ,  �� ��  �� �^  �� �^  �� ��  �� ��      F  , ,  �� v�  �� w�  �� w�  �� v�  �� v�      F  , ,  �� ��  �� �^  �� �^  �� ��  �� ��      F  , ,  �K �&  �K ��  � ��  � �&  �K �&      F  , ,  �� ~�  �� n  �� n  �� ~�  �� ~�      F  , ,  �� ��  �� ��  �� ��  �� ��  �� ��      F  , ,  �K }  �K }�  � }�  � }  �K }      F  , ,  �+ ��  �+ �^  �� �^  �� ��  �+ ��      F  , ,  �K ��  �K �^  � �^  � ��  �K ��      F  , ,  �+ }  �+ }�  �� }�  �� }  �+ }      F  , ,  �K �  �K ��  � ��  � �  �K �      F  , ,  �+ ��  �+ �~  �� �~  �� ��  �+ ��      F  , ,  �K e�  �K fn  � fn  � e�  �K e�      F  , ,  �� d  �� d�  �� d�  �� d  �� d      F  , ,  �� r&  �� r�  �� r�  �� r&  �� r&      F  , ,  �K h�  �K i�  � i�  � h�  �K h�      F  , ,  �+ _f  �+ `.  �� `.  �� _f  �+ _f      F  , ,  �� uF  �� v  �� v  �� uF  �� uF      F  , ,  �� k�  �� l�  �� l�  �� k�  �� k�      F  , ,  �+ b�  �+ cN  �� cN  �� b�  �+ b�      F  , ,  �� jV  �� k  �� k  �� jV  �� jV      F  , ,  �� _f  �� `.  �� `.  �� _f  �� _f      F  , ,  �+ uF  �+ v  �� v  �� uF  �+ uF      F  , ,  �� p�  �� q^  �� q^  �� p�  �� p�      F  , ,  �K mv  �K n>  � n>  � mv  �K mv      F  , ,  �+ d  �+ d�  �� d�  �� d  �+ d      F  , ,  �+ h�  �+ i�  �� i�  �� h�  �+ h�      F  , ,  �� g6  �� g�  �� g�  �� g6  �� g6      F  , ,  �+ o  �+ o�  �� o�  �� o  �+ o      F  , ,  �K `�  �K a�  � a�  � `�  �K `�      F  , ,  �� o  �� o�  �� o�  �� o  �� o      F  , ,  �� _f  �� `.  �� `.  �� _f  �� _f      F  , ,  �+ k�  �+ l�  �� l�  �� k�  �+ k�      F  , ,  �� o  �� o�  �� o�  �� o  �� o      F  , ,  �K \F  �K ]  � ]  � \F  �K \F      F  , ,  �+ jV  �+ k  �� k  �� jV  �+ jV      F  , ,  �� p�  �� q^  �� q^  �� p�  �� p�      F  , ,  �� mv  �� n>  �� n>  �� mv  �� mv      F  , ,  �+ e�  �+ fn  �� fn  �� e�  �+ e�      F  , ,  �+ s�  �+ t~  �� t~  �� s�  �+ s�      F  , ,  �� `�  �� a�  �� a�  �� `�  �� `�      F  , ,  �+ `�  �+ a�  �� a�  �� `�  �+ `�      F  , ,  �K p�  �K q^  � q^  � p�  �K p�      F  , ,  �+ ]�  �+ ^�  �� ^�  �� ]�  �+ ]�      F  , ,  �� k�  �� l�  �� l�  �� k�  �� k�      F  , ,  �� ]�  �� ^�  �� ^�  �� ]�  �� ]�      F  , ,  �+ mv  �+ n>  �� n>  �� mv  �+ mv      F  , ,  �K b�  �K cN  � cN  � b�  �K b�      F  , ,  �� uF  �� v  �� v  �� uF  �� uF      F  , ,  �K g6  �K g�  � g�  � g6  �K g6      F  , ,  �+ g6  �+ g�  �� g�  �� g6  �+ g6      F  , ,  �� e�  �� fn  �� fn  �� e�  �� e�      F  , ,  �� b�  �� cN  �� cN  �� b�  �� b�      F  , ,  �� jV  �� k  �� k  �� jV  �� jV      F  , ,  �K jV  �K k  � k  � jV  �K jV      F  , ,  �� h�  �� i�  �� i�  �� h�  �� h�      F  , ,  �+ \F  �+ ]  �� ]  �� \F  �+ \F      F  , ,  �� b�  �� cN  �� cN  �� b�  �� b�      F  , ,  �+ r&  �+ r�  �� r�  �� r&  �+ r&      F  , ,  �� `�  �� a�  �� a�  �� `�  �� `�      F  , ,  �� h�  �� i�  �� i�  �� h�  �� h�      F  , ,  �� ]�  �� ^�  �� ^�  �� ]�  �� ]�      F  , ,  �K ]�  �K ^�  � ^�  � ]�  �K ]�      F  , ,  �K _f  �K `.  � `.  � _f  �K _f      F  , ,  �K d  �K d�  � d�  � d  �K d      F  , ,  �� s�  �� t~  �� t~  �� s�  �� s�      F  , ,  �� \F  �� ]  �� ]  �� \F  �� \F      F  , ,  �� g6  �� g�  �� g�  �� g6  �� g6      F  , ,  �K o  �K o�  � o�  � o  �K o      F  , ,  �� \F  �� ]  �� ]  �� \F  �� \F      F  , ,  �K k�  �K l�  � l�  � k�  �K k�      F  , ,  �� mv  �� n>  �� n>  �� mv  �� mv      F  , ,  �K uF  �K v  � v  � uF  �K uF      F  , ,  �� r&  �� r�  �� r�  �� r&  �� r&      F  , ,  �K s�  �K t~  � t~  � s�  �K s�      F  , ,  �� e�  �� fn  �� fn  �� e�  �� e�      F  , ,  �� s�  �� t~  �� t~  �� s�  �� s�      F  , ,  �K r&  �K r�  � r�  � r&  �K r&      F  , ,  �+ p�  �+ q^  �� q^  �� p�  �+ p�      F  , ,  �� d  �� d�  �� d�  �� d  �� d      F  , ,  �K @&  �K @�  � @�  � @&  �K @&      F  , ,  �� @&  �� @�  �� @�  �� @&  �� @&      F  , ,  �� @&  �� @�  �� @�  �� @&  �� @&      F  , ,  �+ @&  �+ @�  �� @�  �� @&  �+ @&      F  , ,  �K N6  �K N�  � N�  � N6  �K N6      F  , ,  �+ Y&  �+ Y�  �� Y�  �� Y&  �+ Y&      F  , ,  �� A�  �� B~  �� B~  �� A�  �� A�      F  , ,  �� K  �� K�  �� K�  �� K  �� K      F  , ,  �+ W�  �+ X^  �� X^  �� W�  �+ W�      F  , ,  �� A�  �� B~  �� B~  �� A�  �� A�      F  , ,  �� QV  �� R  �� R  �� QV  �� QV      F  , ,  �K G�  �K H�  � H�  � G�  �K G�      F  , ,  �+ V  �+ V�  �� V�  �� V  �+ V      F  , ,  �� W�  �� X^  �� X^  �� W�  �� W�      F  , ,  �� Ff  �� G.  �� G.  �� Ff  �� Ff      F  , ,  �� I�  �� JN  �� JN  �� I�  �� I�      F  , ,  �+ Tv  �+ U>  �� U>  �� Tv  �+ Tv      F  , ,  �� O�  �� P�  �� P�  �� O�  �� O�      F  , ,  �+ A�  �+ B~  �� B~  �� A�  �+ A�      F  , ,  �K I�  �K JN  � JN  � I�  �K I�      F  , ,  �� Tv  �� U>  �� U>  �� Tv  �� Tv      F  , ,  �+ R�  �+ S�  �� S�  �� R�  �+ R�      F  , ,  �� CF  �� D  �� D  �� CF  �� CF      F  , ,  �K Y&  �K Y�  � Y�  � Y&  �K Y&      F  , ,  �K Ff  �K G.  � G.  � Ff  �K Ff      F  , ,  �� O�  �� P�  �� P�  �� O�  �� O�      F  , ,  �K QV  �K R  � R  � QV  �K QV      F  , ,  �K O�  �K P�  � P�  � O�  �K O�      F  , ,  �K L�  �K Mn  � Mn  � L�  �K L�      F  , ,  �+ QV  �+ R  �� R  �� QV  �+ QV      F  , ,  �� N6  �� N�  �� N�  �� N6  �� N6      F  , ,  �� Y&  �� Y�  �� Y�  �� Y&  �� Y&      F  , ,  �+ O�  �+ P�  �� P�  �� O�  �+ O�      F  , ,  �K W�  �K X^  � X^  � W�  �K W�      F  , ,  �� K  �� K�  �� K�  �� K  �� K      F  , ,  �+ N6  �+ N�  �� N�  �� N6  �+ N6      F  , ,  �K D�  �K E�  � E�  � D�  �K D�      F  , ,  �� D�  �� E�  �� E�  �� D�  �� D�      F  , ,  �� Y&  �� Y�  �� Y�  �� Y&  �� Y&      F  , ,  �+ L�  �+ Mn  �� Mn  �� L�  �+ L�      F  , ,  �� Ff  �� G.  �� G.  �� Ff  �� Ff      F  , ,  �K V  �K V�  � V�  � V  �K V      F  , ,  �+ K  �+ K�  �� K�  �� K  �+ K      F  , ,  �� W�  �� X^  �� X^  �� W�  �� W�      F  , ,  �� G�  �� H�  �� H�  �� G�  �� G�      F  , ,  �K K  �K K�  � K�  � K  �K K      F  , ,  �� N6  �� N�  �� N�  �� N6  �� N6      F  , ,  �� D�  �� E�  �� E�  �� D�  �� D�      F  , ,  �+ I�  �+ JN  �� JN  �� I�  �+ I�      F  , ,  �� V  �� V�  �� V�  �� V  �� V      F  , ,  �K CF  �K D  � D  � CF  �K CF      F  , ,  �+ G�  �+ H�  �� H�  �� G�  �+ G�      F  , ,  �� Tv  �� U>  �� U>  �� Tv  �� Tv      F  , ,  �K Tv  �K U>  � U>  � Tv  �K Tv      F  , ,  �� I�  �� JN  �� JN  �� I�  �� I�      F  , ,  �+ Ff  �+ G.  �� G.  �� Ff  �+ Ff      F  , ,  �� V  �� V�  �� V�  �� V  �� V      F  , ,  �� R�  �� S�  �� S�  �� R�  �� R�      F  , ,  �� L�  �� Mn  �� Mn  �� L�  �� L�      F  , ,  �� R�  �� S�  �� S�  �� R�  �� R�      F  , ,  �+ D�  �+ E�  �� E�  �� D�  �+ D�      F  , ,  �� CF  �� D  �� D  �� CF  �� CF      F  , ,  �� G�  �� H�  �� H�  �� G�  �� G�      F  , ,  �+ CF  �+ D  �� D  �� CF  �+ CF      F  , ,  �� QV  �� R  �� R  �� QV  �� QV      F  , ,  �K A�  �K B~  � B~  � A�  �K A�      F  , ,  �� L�  �� Mn  �� Mn  �� L�  �� L�      F  , ,  �K R�  �K S�  � S�  � R�  �K R�      F  , ,  �+ %�  �+ &^  �� &^  �� %�  �+ %�      F  , ,  �� >�  �� ?^  �� ?^  �� >�  �� >�      F  , ,  �+ .�  �+ /�  �� /�  �� .�  �+ .�      F  , ,  �K '&  �K '�  � '�  � '&  �K '&      F  , ,  �� 9�  �� :�  �� :�  �� 9�  �� 9�      F  , ,  �K 6�  �K 7�  � 7�  � 6�  �K 6�      F  , ,  �� 6�  �� 7�  �� 7�  �� 6�  �� 6�      F  , ,  �K +�  �K ,�  � ,�  � +�  �K +�      F  , ,  �� 3�  �� 4n  �� 4n  �� 3�  �� 3�      F  , ,  �� +�  �� ,�  �� ,�  �� +�  �� +�      F  , ,  �+ +�  �+ ,�  �� ,�  �� +�  �+ +�      F  , ,  �+ 6�  �+ 7�  �� 7�  �� 6�  �+ 6�      F  , ,  �� ;v  �� <>  �� <>  �� ;v  �� ;v      F  , ,  �� (�  �� )~  �� )~  �� (�  �� (�      F  , ,  �� ;v  �� <>  �� <>  �� ;v  �� ;v      F  , ,  �� >�  �� ?^  �� ?^  �� >�  �� >�      F  , ,  �� (�  �� )~  �� )~  �� (�  �� (�      F  , ,  �K 56  �K 5�  � 5�  � 56  �K 56      F  , ,  �+ '&  �+ '�  �� '�  �� '&  �+ '&      F  , ,  �K ;v  �K <>  � <>  � ;v  �K ;v      F  , ,  �� 6�  �� 7�  �� 7�  �� 6�  �� 6�      F  , ,  �+ 3�  �+ 4n  �� 4n  �� 3�  �+ 3�      F  , ,  �K >�  �K ?^  � ?^  � >�  �K >�      F  , ,  �� %�  �� &^  �� &^  �� %�  �� %�      F  , ,  �+ -f  �+ ..  �� ..  �� -f  �+ -f      F  , ,  �+ 0�  �+ 1N  �� 1N  �� 0�  �+ 0�      F  , ,  �+ 8V  �+ 9  �� 9  �� 8V  �+ 8V      F  , ,  �� .�  �� /�  �� /�  �� .�  �� .�      F  , ,  �� *F  �� +  �� +  �� *F  �� *F      F  , ,  �K 3�  �K 4n  � 4n  � 3�  �K 3�      F  , ,  �K *F  �K +  � +  � *F  �K *F      F  , ,  �� 8V  �� 9  �� 9  �� 8V  �� 8V      F  , ,  �� -f  �� ..  �� ..  �� -f  �� -f      F  , ,  �+ >�  �+ ?^  �� ?^  �� >�  �+ >�      F  , ,  �� 2  �� 2�  �� 2�  �� 2  �� 2      F  , ,  �+ =  �+ =�  �� =�  �� =  �+ =      F  , ,  �+ ;v  �+ <>  �� <>  �� ;v  �+ ;v      F  , ,  �K 2  �K 2�  � 2�  � 2  �K 2      F  , ,  �K %�  �K &^  � &^  � %�  �K %�      F  , ,  �� =  �� =�  �� =�  �� =  �� =      F  , ,  �� 56  �� 5�  �� 5�  �� 56  �� 56      F  , ,  �� 0�  �� 1N  �� 1N  �� 0�  �� 0�      F  , ,  �+ 9�  �+ :�  �� :�  �� 9�  �+ 9�      F  , ,  �+ 56  �+ 5�  �� 5�  �� 56  �+ 56      F  , ,  �� '&  �� '�  �� '�  �� '&  �� '&      F  , ,  �+ *F  �+ +  �� +  �� *F  �+ *F      F  , ,  �� .�  �� /�  �� /�  �� .�  �� .�      F  , ,  �� 8V  �� 9  �� 9  �� 8V  �� 8V      F  , ,  �K 9�  �K :�  � :�  � 9�  �K 9�      F  , ,  �� 9�  �� :�  �� :�  �� 9�  �� 9�      F  , ,  �K 0�  �K 1N  � 1N  � 0�  �K 0�      F  , ,  �� 56  �� 5�  �� 5�  �� 56  �� 56      F  , ,  �� *F  �� +  �� +  �� *F  �� *F      F  , ,  �K -f  �K ..  � ..  � -f  �K -f      F  , ,  �� =  �� =�  �� =�  �� =  �� =      F  , ,  �K =  �K =�  � =�  � =  �K =      F  , ,  �+ 2  �+ 2�  �� 2�  �� 2  �+ 2      F  , ,  �K .�  �K /�  � /�  � .�  �K .�      F  , ,  �K (�  �K )~  � )~  � (�  �K (�      F  , ,  �� -f  �� ..  �� ..  �� -f  �� -f      F  , ,  �� 2  �� 2�  �� 2�  �� 2  �� 2      F  , ,  �K 8V  �K 9  � 9  � 8V  �K 8V      F  , ,  �� 0�  �� 1N  �� 1N  �� 0�  �� 0�      F  , ,  �� +�  �� ,�  �� ,�  �� +�  �� +�      F  , ,  �� '&  �� '�  �� '�  �� '&  �� '&      F  , ,  �+ (�  �+ )~  �� )~  �� (�  �+ (�      F  , ,  �� 3�  �� 4n  �� 4n  �� 3�  �� 3�      F  , ,  �� %�  �� &^  �� &^  �� %�  �� %�      F  , ,  �� 	v  �� 
>  �� 
>  �� 	v  �� 	v      F  , ,  �K 	v  �K 
>  � 
>  � 	v  �K 	v      F  , ,  �+ 	v  �+ 
>  �� 
>  �� 	v  �+ 	v      F  , ,  �� 	v  �� 
>  �� 
>  �� 	v  �� 	v      F  , ,  �K f  �K .  � .  � f  �K f      F  , ,  �� "v  �� #>  �� #>  �� "v  �� "v      F  , ,  �K 6  �K �  � �  � 6  �K 6      F  , ,  �� �  �� ~  �� ~  �� �  �� �      F  , ,  �+ �  �+ ^  �� ^  �� �  �+ �      F  , ,  �+ F  �+   ��   �� F  �+ F      F  , ,  �+   �+ �  �� �  ��   �+       F  , ,  �� f  �� .  �� .  �� f  �� f      F  , ,  �� �  �� N  �� N  �� �  �� �      F  , ,  �K �  �K ^  � ^  � �  �K �      F  , ,  �+ �  �+ N  �� N  �� �  �+ �      F  , ,  �K  �  �K !�  � !�  �  �  �K  �      F  , ,  �K "v  �K #>  � #>  � "v  �K "v      F  , ,  �K   �K �  � �  �   �K       F  , ,  �� 6  �� �  �� �  �� 6  �� 6      F  , ,  �+ �  �+ �  �� �  �� �  �+ �      F  , ,  ��   �� �  �� �  ��   ��       F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �� 6  �� �  �� �  �� 6  �� 6      F  , ,  �+ f  �+ .  �� .  �� f  �+ f      F  , ,  ��   �� �  �� �  ��   ��       F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �� &  �� �  �� �  �� &  �� &      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �� F  ��   ��   �� F  �� F      F  , ,  ��  �  �� !�  �� !�  ��  �  ��  �      F  , ,  ��  �  �� !�  �� !�  ��  �  ��  �      F  , ,  �� F  ��   ��   �� F  �� F      F  , ,  �� $  �� $�  �� $�  �� $  �� $      F  , ,  �K   �K �  � �  �   �K       F  , ,  �+ �  �+ n  �� n  �� �  �+ �      F  , ,  �+ �  �+ ~  �� ~  �� �  �+ �      F  , ,  �K &  �K �  � �  � &  �K &      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �+ $  �+ $�  �� $�  �� $  �+ $      F  , ,  �� �  �� ~  �� ~  �� �  �� �      F  , ,  �+ "v  �+ #>  �� #>  �� "v  �+ "v      F  , ,  ��   �� �  �� �  ��   ��       F  , ,  �K �  �K �  � �  � �  �K �      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �� �  �� N  �� N  �� �  �� �      F  , ,  �K �  �K N  � N  � �  �K �      F  , ,  �+ �  �+ �  �� �  �� �  �+ �      F  , ,  �K �  �K n  � n  � �  �K �      F  , ,  �+  �  �+ !�  �� !�  ��  �  �+  �      F  , ,  �� V  ��    ��    �� V  �� V      F  , ,  �� &  �� �  �� �  �� &  �� &      F  , ,  �K F  �K   �   � F  �K F      F  , ,  �� �  �� ^  �� ^  �� �  �� �      F  , ,  �K V  �K    �    � V  �K V      F  , ,  �� "v  �� #>  �� #>  �� "v  �� "v      F  , ,  �+ V  �+    ��    �� V  �+ V      F  , ,  �� V  ��    ��    �� V  �� V      F  , ,  �+ &  �+ �  �� �  �� &  �+ &      F  , ,  �� �  �� ^  �� ^  �� �  �� �      F  , ,  �� $  �� $�  �� $�  �� $  �� $      F  , ,  �K �  �K �  � �  � �  �K �      F  , ,  �K �  �K �  � �  � �  �K �      F  , ,  �K �  �K ~  � ~  � �  �K �      F  , ,  �+ �  �+ �  �� �  �� �  �+ �      F  , ,  �� �  �� n  �� n  �� �  �� �      F  , ,  �� f  �� .  �� .  �� f  �� f      F  , ,  �+ 6  �+ �  �� �  �� 6  �+ 6      F  , ,  �K $  �K $�  � $�  � $  �K $      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �+   �+ �  �� �  ��   �+       F  , ,  ��   �� �  �� �  ��   ��       F  , ,  �� �  �� n  �� n  �� �  �� �      F  , ,  ��  �  ��  �^  ��  �^  ��  �  ��  �      F  , ,  �+  ��  �+  ��  ��  ��  ��  ��  �+  ��      F  , ,  ��  ��  ��  �~  ��  �~  ��  ��  ��  ��      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  ��  ��  ��  �N  ��  �N  ��  ��  ��  ��      F  , ,  �K  ��  �K  ��  �  ��  �  ��  �K  ��      F  , ,  �+  ��  �+  �~  ��  �~  ��  ��  �+  ��      F  , ,  �K �  �K �  � �  � �  �K �      F  , ,  ��  �F  ��  �  ��  �  ��  �F  ��  �F      F  , ,  ��  �v  ��  �>  ��  �>  ��  �v  ��  �v      F  , ,  ��  �f  ��  �.  ��  �.  ��  �f  ��  �f      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �K  �F  �K  �  �  �  �  �F  �K  �F      F  , ,  �K  �f  �K  �.  �  �.  �  �f  �K  �f      F  , ,  �+  �&  �+  ��  ��  ��  ��  �&  �+  �&      F  , ,  ��    ��  �  ��  �  ��    ��        F  , ,  �� V  ��   ��   �� V  �� V      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �� �  �� �  �� �  �� �  �� �      F  , ,  �+  �  �+  ��  ��  ��  ��  �  �+  �      F  , ,  �+ �  �+ n  �� n  �� �  �+ �      F  , ,  �+ �  �+ �  �� �  �� �  �+ �      F  , ,  �K  ��  �K  �  �  �  �  ��  �K  ��      F  , ,  ��  ��  ��  �~  ��  �~  ��  ��  ��  ��      F  , ,  ��  �v  ��  �>  ��  �>  ��  �v  ��  �v      F  , ,  �+ 6  �+ �  �� �  �� 6  �+ 6      F  , ,  �+ V  �+   ��   �� V  �+ V      F  , ,  ��  �F  ��  �  ��  �  ��  �F  ��  �F      F  , ,  �+  ��  �+  �N  ��  �N  ��  ��  �+  ��      F  , ,  ��  �  ��  �^  ��  �^  ��  �  ��  �      F  , ,  �K  �v  �K  �>  �  �>  �  �v  �K  �v      F  , ,  �� 6  �� �  �� �  �� 6  �� 6      F  , ,  ��  ��  ��  �  ��  �  ��  ��  ��  ��      F  , ,  �+  ��  �+  ��  ��  ��  ��  ��  �+  ��      F  , ,  �K �  �K �  � �  � �  �K �      F  , ,  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��      F  , ,  ��  �  ��  ��  ��  ��  ��  �  ��  �      F  , ,  �+  ��  �+  �  ��  �  ��  ��  �+  ��      F  , ,  ��  �  ��  ��  ��  ��  ��  �  ��  �      F  , ,  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��      F  , ,  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��      F  , ,  ��  �&  ��  ��  ��  ��  ��  �&  ��  �&      F  , ,  �� 6  �� �  �� �  �� 6  �� 6      F  , ,  �K  �  �K  ��  �  ��  �  �  �K  �      F  , ,  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��      F  , ,  �+ �  �+ �  �� �  �� �  �+ �      F  , ,  �K  �&  �K  ��  �  ��  �  �&  �K  �&      F  , ,  �K �  �K n  � n  � �  �K �      F  , ,  �K V  �K   �   � V  �K V      F  , ,  �K    �K  �  �  �  �    �K        F  , ,  ��  ��  ��  �N  ��  �N  ��  ��  ��  ��      F  , ,  �� �  �� n  �� n  �� �  �� �      F  , ,  �+  �F  �+  �  ��  �  ��  �F  �+  �F      F  , ,  �� V  ��   ��   �� V  �� V      F  , ,  ��  �&  ��  ��  ��  ��  ��  �&  ��  �&      F  , ,  ��    ��  �  ��  �  ��    ��        F  , ,  �K  �  �K  �^  �  �^  �  �  �K  �      F  , ,  ��  �f  ��  �.  ��  �.  ��  �f  ��  �f      F  , ,  �+  �  �+  �^  ��  �^  ��  �  �+  �      F  , ,  �K 6  �K �  � �  � 6  �K 6      F  , ,  �K  ��  �K  �N  �  �N  �  ��  �K  ��      F  , ,  �+    �+  �  ��  �  ��    �+        F  , ,  �+  �v  �+  �>  ��  �>  ��  �v  �+  �v      F  , ,  �K  ��  �K  ��  �  ��  �  ��  �K  ��      F  , ,  ��  ��  ��  �  ��  �  ��  ��  ��  ��      F  , ,  �+  �f  �+  �.  ��  �.  ��  �f  �+  �f      F  , ,  �� �  �� n  �� n  �� �  �� �      F  , ,  �K  ��  �K  �~  �  �~  �  ��  �K  ��      F  , , 
s Z� 
s [~ ; [~ ; Z� 
s Z�      F  , , � Z� � [~ [ [~ [ Z� � Z�      F  , ,  Z�  [~ � [~ � Z�  Z�      F  , , � Z� � [~ 	� [~ 	� Z� � Z�      F  , , � �f � �. [ �. [ �f � �f      F  , ,  �f  �. � �. � �f  �f      F  , , � �f � �. 	� �. 	� �f � �f      F  , , 
s �f 
s �. ; �. ; �f 
s �f      F  , , � �� � �� [ �� [ �� � ��      F  , , � �� � �� 	� �� 	� �� � ��      F  , ,  ��  �� � �� � ��  ��      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , , 
s � 
s �� ; �� ; � 
s �      F  , ,  ��  �� � �� � ��  ��      F  , ,  ��  �N � �N � ��  ��      F  , ,  �  �� � �� � �  �      F  , , 
s �� 
s �^ ; �^ ; �� 
s ��      F  , ,  ��  �n � �n � ��  ��      F  , ,  �V  � � � � �V  �V      F  , , 
s �f 
s �. ; �. ; �f 
s �f      F  , ,  �6  �� � �� � �6  �6      F  , , � �� � ž 	� ž 	� �� � ��      F  , , 
s �v 
s �> ; �> ; �v 
s �v      F  , , � Ɔ � �N 	� �N 	� Ɔ � Ɔ      F  , , 
s �� 
s  ;  ; �� 
s ��      F  , , � �f � �. 	� �. 	� �f � �f      F  , ,  Ɔ  �N � �N � Ɔ  Ɔ      F  , , � Ɔ � �N [ �N [ Ɔ � Ɔ      F  , ,  ��  ž � ž � ��  ��      F  , , 
s �& 
s �� ; �� ; �& 
s �&      F  , , 
s �� 
s �N ; �N ; �� 
s ��      F  , ,  ��  �� � �� � ��  ��      F  , , � �� � �N [ �N [ �� � ��      F  , , 
s �� 
s �n ; �n ; �� 
s ��      F  , , � � � �� [ �� [ � � �      F  , , 
s Ɔ 
s �N ; �N ; Ɔ 
s Ɔ      F  , ,  �v  �> � �> � �v  �v      F  , , � �� � �n [ �n [ �� � ��      F  , , 
s � 
s �� ; �� ; � 
s �      F  , , 
s �� 
s �~ ; �~ ; �� 
s ��      F  , , � �� � �N 	� �N 	� �� � ��      F  , , � �6 � �� [ �� [ �6 � �6      F  , , 
s �6 
s �� ; �� ; �6 
s �6      F  , , � � � �� 	� �� 	� � � �      F  , , � �� � �� [ �� [ �� � ��      F  , ,  �  �� � �� � �  �      F  , , � �� � �n 	� �n 	� �� � ��      F  , , � �V � � [ � [ �V � �V      F  , , � �6 � �� 	� �� 	� �6 � �6      F  , , � �� � �� [ �� [ �� � ��      F  , , � �� � �� 	� �� 	� �� � ��      F  , ,  ��  �^ � �^ � ��  ��      F  , , � �v � �> [ �> [ �v � �v      F  , , � �V � � 	� � 	� �V � �V      F  , , � � � �� [ �� [ � � �      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , ,  �&  �� � �� � �&  �&      F  , , 
s �� 
s ž ; ž ; �� 
s ��      F  , , � �� � �� 	� �� 	� �� � ��      F  , , � �� � �^ [ �^ [ �� � ��      F  , , � �v � �> 	� �> 	� �v � �v      F  , , � �& � �� [ �� [ �& � �&      F  , ,  ��  �~ � �~ � ��  ��      F  , , � � � �� 	� �� 	� � � �      F  , , 
s �F 
s � ; � ; �F 
s �F      F  , , � �� � �~ [ �~ [ �� � ��      F  , ,  �F  � � � � �F  �F      F  , , 
s �V 
s � ; � ; �V 
s �V      F  , , � �� � �^ 	� �^ 	� �� � ��      F  , , � �F � � [ � [ �F � �F      F  , , � �& � �� 	� �� 	� �& � �&      F  , , � �� �  [  [ �� � ��      F  , ,  ��   �  � ��  ��      F  , , � �� � �~ 	� �~ 	� �� � ��      F  , , � �f � �. [ �. [ �f � �f      F  , ,  �f  �. � �. � �f  �f      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , , � �F � � 	� � 	� �F � �F      F  , , � �� � ž [ ž [ �� � ��      F  , , � �� �  	�  	� �� � ��      F  , ,  �  �� � �� � �  �      F  , , � �� � �� [ �� [ �� � ��      F  , , 
s �V 
s � ; � ; �V 
s �V      F  , , 
s �� 
s �n ; �n ; �� 
s ��      F  , ,  �F  � � � � �F  �F      F  , , � �� � �~ 	� �~ 	� �� � ��      F  , ,  �&  �� � �� � �&  �&      F  , ,  ��  �� � �� � ��  ��      F  , , � �& � �� [ �� [ �& � �&      F  , , 
s �F 
s � ; � ; �F 
s �F      F  , ,  ��  �� � �� � ��  ��      F  , , � �f � �. [ �. [ �f � �f      F  , , 
s �f 
s �. ; �. ; �f 
s �f      F  , , � �F � � [ � [ �F � �F      F  , , � �� � �N [ �N [ �� � ��      F  , , � �V � � [ � [ �V � �V      F  , ,  ��  �~ � �~ � ��  ��      F  , , 
s �� 
s �~ ; �~ ; �� 
s ��      F  , , � �� � �� 	� �� 	� �� � ��      F  , , � �� � �� 	� �� 	� �� � ��      F  , , � �V � � 	� � 	� �V � �V      F  , ,  ��  �N � �N � ��  ��      F  , ,  �6  �� � �� � �6  �6      F  , , � �v � �> [ �> [ �v � �v      F  , , � � � �� [ �� [ � � �      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , , 
s �� 
s �N ; �N ; �� 
s ��      F  , ,  �v  �> � �> � �v  �v      F  , , � �� � �� [ �� [ �� � ��      F  , , � �� � �� [ �� [ �� � ��      F  , , � �� � �n [ �n [ �� � ��      F  , , � �v � �> 	� �> 	� �v � �v      F  , , 
s �v 
s �> ; �> ; �v 
s �v      F  , , � �� � �n 	� �n 	� �� � ��      F  , , � �� � �� 	� �� 	� �� � ��      F  , , 
s � 
s �� ; �� ; � 
s �      F  , ,  �V  � � � � �V  �V      F  , , � �6 � �� [ �� [ �6 � �6      F  , ,  �  �� � �� � �  �      F  , , � � � �� 	� �� 	� � � �      F  , , 
s �& 
s �� ; �� ; �& 
s �&      F  , , � � � �� [ �� [ � � �      F  , , 
s �6 
s �� ; �� ; �6 
s �6      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , , � � � �� 	� �� 	� � � �      F  , , � �& � �� 	� �� 	� �& � �&      F  , , 
s �� 
s �^ ; �^ ; �� 
s ��      F  , , � �f � �. 	� �. 	� �f � �f      F  , , � �� � �~ [ �~ [ �� � ��      F  , ,  ��  �^ � �^ � ��  ��      F  , , � �� � �� 	� �� 	� �� � ��      F  , , � �6 � �� 	� �� 	� �6 � �6      F  , ,  �f  �. � �. � �f  �f      F  , , 
s � 
s �� ; �� ; � 
s �      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , ,  ��  �n � �n � ��  ��      F  , , � �� � �^ [ �^ [ �� � ��      F  , ,  ��  �� � �� � ��  ��      F  , , � �� � �N 	� �N 	� �� � ��      F  , , � �F � � 	� � 	� �F � �F      F  , ,  ��  �� � �� � ��  ��      F  , , � �� � �� [ �� [ �� � ��      F  , , � �� � �^ 	� �^ 	� �� � ��      F  , , � �� � �� 	� �� 	� �� � ��      F  , , 
s �F 
s � ; � ; �F 
s �F      F  , , � y� � z� 	� z� 	� y� � y�      F  , , 
s } 
s }� ; }� ; } 
s }      F  , , � {� � |N 	� |N 	� {� � {�      F  , , 
s xf 
s y. ; y. ; xf 
s xf      F  , ,  {�  |N � |N � {�  {�      F  , , 
s � 
s �� ; �� ; � 
s �      F  , , � �� � �~ 	� �~ 	� �� � ��      F  , ,  �  �� � �� � �  �      F  , ,  xf  y. � y. � xf  xf      F  , , � } � }� 	� }� 	� } � }      F  , ,  ��  �^ � �^ � ��  ��      F  , , � �� � �^ 	� �^ 	� �� � ��      F  , ,  }  }� � }� � }  }      F  , , � �� � �� [ �� [ �� � ��      F  , , 
s ~� 
s n ; n ; ~� 
s ~�      F  , , � �V � � 	� � 	� �V � �V      F  , ,  �&  �� � �� � �&  �&      F  , , � �� � �^ [ �^ [ �� � ��      F  , , � ~� � n [ n [ ~� � ~�      F  , , � v� � w� [ w� [ v� � v�      F  , , 
s �� 
s �^ ; �^ ; �� 
s ��      F  , , � �F � � 	� � 	� �F � �F      F  , , � �v � �> [ �> [ �v � �v      F  , ,  ��  �~ � �~ � ��  ��      F  , , � �� � �� [ �� [ �� � ��      F  , , � �& � �� 	� �� 	� �& � �&      F  , , 
s �6 
s �� ; �� ; �6 
s �6      F  , ,  �F  � � � � �F  �F      F  , , � ~� � n 	� n 	� ~� � ~�      F  , , 
s y� 
s z� ; z� ; y� 
s y�      F  , , � �F � � [ � [ �F � �F      F  , , 
s {� 
s |N ; |N ; {� 
s {�      F  , ,  ��  �� � �� � ��  ��      F  , , � �V � � [ � [ �V � �V      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , , � xf � y. [ y. [ xf � xf      F  , , 
s �v 
s �> ; �> ; �v 
s �v      F  , , � �v � �> 	� �> 	� �v � �v      F  , ,  �V  � � � � �V  �V      F  , , 
s �& 
s �� ; �� ; �& 
s �&      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , , � �& � �� [ �� [ �& � �&      F  , ,  ��  �� � �� � ��  ��      F  , , � �� � �� 	� �� 	� �� � ��      F  , , � �� � �� 	� �� 	� �� � ��      F  , ,  �6  �� � �� � �6  �6      F  , , 
s �� 
s �� ; �� ; �� 
s ��      F  , ,  y�  z� � z� � y�  y�      F  , , � y� � z� [ z� [ y� � y�      F  , , � �� � �~ [ �~ [ �� � ��      F  , , � �6 � �� 	� �� 	� �6 � �6      F  , ,  ��  �� � �� � ��  ��      F  , , � �� � �� [ �� [ �� � ��      F  , ,  v�  w� � w� � v�  v�      F  , ,  �v  �> � �> � �v  �v      F  , , � v� � w� 	� w� 	� v� � v�      F  , , � �6 � �� [ �� [ �6 � �6      F  , , � {� � |N [ |N [ {� � {�      F  , , 
s �V 
s � ; � ; �V 
s �V      F  , ,  ~�  n � n � ~�  ~�      F  , , 
s �� 
s �~ ; �~ ; �� 
s ��      F  , , � � � �� 	� �� 	� � � �      F  , , � � � �� [ �� [ � � �      F  , , � xf � y. 	� y. 	� xf � xf      F  , , 
s v� 
s w� ; w� ; v� 
s v�      F  , , � } � }� [ }� [ } � }      F  , , � g6 � g� 	� g� 	� g6 � g6      F  , ,  `�  a� � a� � `�  `�      F  , , � `� � a� 	� a� 	� `� � `�      F  , , � _f � `. [ `. [ _f � _f      F  , , 
s s� 
s t~ ; t~ ; s� 
s s�      F  , , � jV � k [ k [ jV � jV      F  , , � `� � a� [ a� [ `� � `�      F  , ,  _f  `. � `. � _f  _f      F  , , 
s `� 
s a� ; a� ; `� 
s `�      F  , ,  g6  g� � g� � g6  g6      F  , , � b� � cN 	� cN 	� b� � b�      F  , , � d � d� [ d� [ d � d      F  , ,  k�  l� � l� � k�  k�      F  , , � s� � t~ 	� t~ 	� s� � s�      F  , , � k� � l� [ l� [ k� � k�      F  , , 
s uF 
s v ; v ; uF 
s uF      F  , ,  s�  t~ � t~ � s�  s�      F  , , � uF � v [ v [ uF � uF      F  , , � o � o� 	� o� 	� o � o      F  , , � _f � `. 	� `. 	� _f � _f      F  , , � e� � fn 	� fn 	� e� � e�      F  , ,  b�  cN � cN � b�  b�      F  , , � r& � r� 	� r� 	� r& � r&      F  , , � mv � n> [ n> [ mv � mv      F  , ,  h�  i� � i� � h�  h�      F  , ,  ]�  ^� � ^� � ]�  ]�      F  , , 
s mv 
s n> ; n> ; mv 
s mv      F  , , 
s r& 
s r� ; r� ; r& 
s r&      F  , , � mv � n> 	� n> 	� mv � mv      F  , , 
s jV 
s k ; k ; jV 
s jV      F  , , 
s d 
s d� ; d� ; d 
s d      F  , , � p� � q^ [ q^ [ p� � p�      F  , , 
s \F 
s ] ; ] ; \F 
s \F      F  , , 
s g6 
s g� ; g� ; g6 
s g6      F  , ,  e�  fn � fn � e�  e�      F  , , � ]� � ^� [ ^� [ ]� � ]�      F  , , 
s ]� 
s ^� ; ^� ; ]� 
s ]�      F  , , � g6 � g� [ g� [ g6 � g6      F  , , 
s b� 
s cN ; cN ; b� 
s b�      F  , , 
s k� 
s l� ; l� ; k� 
s k�      F  , , � jV � k 	� k 	� jV � jV      F  , , 
s o 
s o� ; o� ; o 
s o      F  , , � h� � i� 	� i� 	� h� � h�      F  , ,  jV  k � k � jV  jV      F  , ,  \F  ] � ] � \F  \F      F  , , � s� � t~ [ t~ [ s� � s�      F  , , � b� � cN [ cN [ b� � b�      F  , ,  uF  v � v � uF  uF      F  , , � r& � r� [ r� [ r& � r&      F  , , � \F � ] 	� ] 	� \F � \F      F  , , � d � d� 	� d� 	� d � d      F  , , � o � o� [ o� [ o � o      F  , , � ]� � ^� 	� ^� 	� ]� � ]�      F  , ,  r&  r� � r� � r&  r&      F  , , 
s h� 
s i� ; i� ; h� 
s h�      F  , ,  mv  n> � n> � mv  mv      F  , , � \F � ] [ ] [ \F � \F      F  , ,  p�  q^ � q^ � p�  p�      F  , , � k� � l� 	� l� 	� k� � k�      F  , ,  d  d� � d� � d  d      F  , , 
s e� 
s fn ; fn ; e� 
s e�      F  , , � e� � fn [ fn [ e� � e�      F  , , 
s p� 
s q^ ; q^ ; p� 
s p�      F  , ,  o  o� � o� � o  o      F  , , � p� � q^ 	� q^ 	� p� � p�      F  , , 
s _f 
s `. ; `. ; _f 
s _f      F  , , � uF � v 	� v 	� uF � uF      F  , , � h� � i� [ i� [ h� � h�      F  , , 
s @& 
s @� ; @� ; @& 
s @&      F  , , � @& � @� 	� @� 	� @& � @&      F  , , � @& � @� [ @� [ @& � @&      F  , ,  @&  @� � @� � @&  @&      F  , , � N6 � N� 	� N� 	� N6 � N6      F  , , � Ff � G. 	� G. 	� Ff � Ff      F  , , 
s K 
s K� ; K� ; K 
s K      F  , ,  W�  X^ � X^ � W�  W�      F  , , 
s V 
s V� ; V� ; V 
s V      F  , , � O� � P� 	� P� 	� O� � O�      F  , , 
s I� 
s JN ; JN ; I� 
s I�      F  , , 
s Y& 
s Y� ; Y� ; Y& 
s Y&      F  , ,  Tv  U> � U> � Tv  Tv      F  , , � N6 � N� [ N� [ N6 � N6      F  , , � G� � H� [ H� [ G� � G�      F  , , � QV � R 	� R 	� QV � QV      F  , , � Tv � U> [ U> [ Tv � Tv      F  , ,  L�  Mn � Mn � L�  L�      F  , ,  O�  P� � P� � O�  O�      F  , ,  QV  R � R � QV  QV      F  , , � G� � H� 	� H� 	� G� � G�      F  , , � L� � Mn [ Mn [ L� � L�      F  , , 
s O� 
s P� ; P� ; O� 
s O�      F  , ,  D�  E� � E� � D�  D�      F  , ,  CF  D � D � CF  CF      F  , ,  Ff  G. � G. � Ff  Ff      F  , , 
s CF 
s D ; D ; CF 
s CF      F  , ,  Y&  Y� � Y� � Y&  Y&      F  , , � V � V� [ V� [ V � V      F  , , � CF � D [ D [ CF � CF      F  , , � R� � S� 	� S� 	� R� � R�      F  , , � I� � JN 	� JN 	� I� � I�      F  , ,  R�  S� � S� � R�  R�      F  , , 
s Tv 
s U> ; U> ; Tv 
s Tv      F  , , � D� � E� [ E� [ D� � D�      F  , ,  I�  JN � JN � I�  I�      F  , , � D� � E� 	� E� 	� D� � D�      F  , , � A� � B~ 	� B~ 	� A� � A�      F  , , 
s N6 
s N� ; N� ; N6 
s N6      F  , ,  A�  B~ � B~ � A�  A�      F  , , � O� � P� [ P� [ O� � O�      F  , ,  K  K� � K� � K  K      F  , , � Tv � U> 	� U> 	� Tv � Tv      F  , , � I� � JN [ JN [ I� � I�      F  , , 
s G� 
s H� ; H� ; G� 
s G�      F  , , � R� � S� [ S� [ R� � R�      F  , , 
s Ff 
s G. ; G. ; Ff 
s Ff      F  , , � W� � X^ [ X^ [ W� � W�      F  , , 
s W� 
s X^ ; X^ ; W� 
s W�      F  , , � V � V� 	� V� 	� V � V      F  , , � K � K� 	� K� 	� K � K      F  , ,  G�  H� � H� � G�  G�      F  , , � CF � D 	� D 	� CF � CF      F  , ,  V  V� � V� � V  V      F  , , � QV � R [ R [ QV � QV      F  , , 
s QV 
s R ; R ; QV 
s QV      F  , , 
s L� 
s Mn ; Mn ; L� 
s L�      F  , , 
s A� 
s B~ ; B~ ; A� 
s A�      F  , , � Ff � G. [ G. [ Ff � Ff      F  , , � W� � X^ 	� X^ 	� W� � W�      F  , ,  N6  N� � N� � N6  N6      F  , , � L� � Mn 	� Mn 	� L� � L�      F  , , � K � K� [ K� [ K � K      F  , , � A� � B~ [ B~ [ A� � A�      F  , , � Y& � Y� [ Y� [ Y& � Y&      F  , , 
s R� 
s S� ; S� ; R� 
s R�      F  , , � Y& � Y� 	� Y� 	� Y& � Y&      F  , , 
s D� 
s E� ; E� ; D� 
s D�      F  , ,  2  2� � 2� � 2  2      F  , , � 3� � 4n [ 4n [ 3� � 3�      F  , , � 6� � 7� 	� 7� 	� 6� � 6�      F  , , � (� � )~ 	� )~ 	� (� � (�      F  , , � 0� � 1N 	� 1N 	� 0� � 0�      F  , , 
s +� 
s ,� ; ,� ; +� 
s +�      F  , , � >� � ?^ [ ?^ [ >� � >�      F  , , � *F � + [ + [ *F � *F      F  , , � 0� � 1N [ 1N [ 0� � 0�      F  , ,  (�  )~ � )~ � (�  (�      F  , ,  0�  1N � 1N � 0�  0�      F  , ,  9�  :� � :� � 9�  9�      F  , , � .� � /� 	� /� 	� .� � .�      F  , , � +� � ,� 	� ,� 	� +� � +�      F  , , � *F � + 	� + 	� *F � *F      F  , , � 56 � 5� 	� 5� 	� 56 � 56      F  , , � -f � .. 	� .. 	� -f � -f      F  , , � 2 � 2� 	� 2� 	� 2 � 2      F  , , � .� � /� [ /� [ .� � .�      F  , , � %� � &^ 	� &^ 	� %� � %�      F  , ,  56  5� � 5� � 56  56      F  , , � +� � ,� [ ,� [ +� � +�      F  , ,  '&  '� � '� � '&  '&      F  , , � ;v � <> [ <> [ ;v � ;v      F  , , � = � =� 	� =� 	� = � =      F  , , 
s 2 
s 2� ; 2� ; 2 
s 2      F  , , � 56 � 5� [ 5� [ 56 � 56      F  , ,  3�  4n � 4n � 3�  3�      F  , ,  8V  9 � 9 � 8V  8V      F  , , 
s 3� 
s 4n ; 4n ; 3� 
s 3�      F  , , 
s %� 
s &^ ; &^ ; %� 
s %�      F  , ,  .�  /� � /� � .�  .�      F  , , � 8V � 9 [ 9 [ 8V � 8V      F  , , 
s >� 
s ?^ ; ?^ ; >� 
s >�      F  , , 
s 8V 
s 9 ; 9 ; 8V 
s 8V      F  , , � 9� � :� [ :� [ 9� � 9�      F  , ,  +�  ,� � ,� � +�  +�      F  , , � '& � '� [ '� [ '& � '&      F  , ,  ;v  <> � <> � ;v  ;v      F  , , � (� � )~ [ )~ [ (� � (�      F  , , � '& � '� 	� '� 	� '& � '&      F  , , � ;v � <> 	� <> 	� ;v � ;v      F  , , 
s = 
s =� ; =� ; = 
s =      F  , ,  >�  ?^ � ?^ � >�  >�      F  , , � %� � &^ [ &^ [ %� � %�      F  , , � 8V � 9 	� 9 	� 8V � 8V      F  , , � 9� � :� 	� :� 	� 9� � 9�      F  , , � 6� � 7� [ 7� [ 6� � 6�      F  , , 
s -f 
s .. ; .. ; -f 
s -f      F  , ,  -f  .. � .. � -f  -f      F  , , 
s *F 
s + ; + ; *F 
s *F      F  , ,  =  =� � =� � =  =      F  , , 
s 56 
s 5� ; 5� ; 56 
s 56      F  , , � -f � .. [ .. [ -f � -f      F  , , 
s (� 
s )~ ; )~ ; (� 
s (�      F  , , � 3� � 4n 	� 4n 	� 3� � 3�      F  , ,  6�  7� � 7� � 6�  6�      F  , , 
s 0� 
s 1N ; 1N ; 0� 
s 0�      F  , , 
s ;v 
s <> ; <> ; ;v 
s ;v      F  , , � >� � ?^ 	� ?^ 	� >� � >�      F  , , � 2 � 2� [ 2� [ 2 � 2      F  , ,  %�  &^ � &^ � %�  %�      F  , , � = � =� [ =� [ = � =      F  , , 
s 6� 
s 7� ; 7� ; 6� 
s 6�      F  , , 
s .� 
s /� ; /� ; .� 
s .�      F  , ,  *F  + � + � *F  *F      F  , , 
s 9� 
s :� ; :� ; 9� 
s 9�      F  , , 
s '& 
s '� ; '� ; '& 
s '&      F  , ,  	v  
> � 
> � 	v  	v      F  , , � 	v � 
> 	� 
> 	� 	v � 	v      F  , , 
s 	v 
s 
> ; 
> ; 	v 
s 	v      F  , , � 	v � 
> [ 
> [ 	v � 	v      F  , , � $ � $� [ $� [ $ � $      F  , , � � � ~ 	� ~ 	� � � �      F  , , � � � ^ [ ^ [ � � �      F  , , � � � n 	� n 	� � � �      F  , , � $ � $� 	� $� 	� $ � $      F  , ,    � � � �         F  , , � � � � 	� � 	� � � �      F  , , 
s $ 
s $� ; $� ; $ 
s $      F  , ,  F   �  � F  F      F  , , � F �  [  [ F � F      F  , , � f � . [ . [ f � f      F  , , 
s  � 
s !� ; !� ;  � 
s  �      F  , , 
s & 
s � ; � ; & 
s &      F  , , �  � � !� [ !� [  � �  �      F  , , 
s � 
s ^ ; ^ ; � 
s �      F  , , 
s F 
s  ;  ; F 
s F      F  , , � V �   [   [ V � V      F  , ,  V    �   � V  V      F  , , � � � � [ � [ � � �      F  , ,  �  ~ � ~ � �  �      F  , , � & � � [ � [ & � &      F  , , �  � � !� 	� !� 	�  � �  �      F  , , � � � � [ � [ � � �      F  , , 
s  
s � ; � ;  
s       F  , , � & � � 	� � 	� & � &      F  , , � f � . 	� . 	� f � f      F  , ,  �  n � n � �  �      F  , , 
s 6 
s � ; � ; 6 
s 6      F  , , � � � � [ � [ � � �      F  , , 
s � 
s � ; � ; � 
s �      F  , ,  $  $� � $� � $  $      F  , , �  � � [ � [  �       F  , , � � � � 	� � 	� � � �      F  , , � � � � 	� � 	� � � �      F  , , � 6 � � 	� � 	� 6 � 6      F  , , � 6 � � [ � [ 6 � 6      F  , , 
s V 
s   ;   ; V 
s V      F  , ,  �  N � N � �  �      F  , ,    � � � �         F  , ,  "v  #> � #> � "v  "v      F  , , 
s � 
s N ; N ; � 
s �      F  , ,  &  � � � � &  &      F  , ,   �  !� � !� �  �   �      F  , ,  �  � � � � �  �      F  , , � V �   	�   	� V � V      F  , , � � � N 	� N 	� � � �      F  , ,  �  ^ � ^ � �  �      F  , , 
s � 
s � ; � ; � 
s �      F  , , � � � n [ n [ � � �      F  , , � � � N [ N [ � � �      F  , , 
s � 
s n ; n ; � 
s �      F  , ,  �  � � � � �  �      F  , , 
s f 
s . ; . ; f 
s f      F  , , �  � � 	� � 	�  �       F  , , �  � � [ � [  �       F  , , � F �  	�  	� F � F      F  , , 
s  
s � ; � ;  
s       F  , , � � � ^ 	� ^ 	� � � �      F  , , � "v � #> [ #> [ "v � "v      F  , , � � � ~ [ ~ [ � � �      F  , , � "v � #> 	� #> 	� "v � "v      F  , , �  � � 	� � 	�  �       F  , ,  6  � � � � 6  6      F  , , 
s "v 
s #> ; #> ; "v 
s "v      F  , , 
s � 
s ~ ; ~ ; � 
s �      F  , ,  �  � � � � �  �      F  , ,  f  . � . � f  f      F  , , 
s � 
s � ; � ; � 
s �      F  , ,   �f   �. �  �. �  �f   �f      F  , , 
s  �� 
s  �~ ;  �~ ;  �� 
s  ��      F  , , � 6 � � 	� � 	� 6 � 6      F  , ,  �  � � � � �  �      F  , , �  �� �  �� 	�  �� 	�  �� �  ��      F  , ,   ��   �� �  �� �  ��   ��      F  , , � � � � 	� � 	� � � �      F  , , �  � �  �^ 	�  �^ 	�  � �  �      F  , , �  �v �  �> 	�  �> 	�  �v �  �v      F  , , �  �� �  � [  � [  �� �  ��      F  , , 
s � 
s � ; � ; � 
s �      F  , , �  �� �  �� 	�  �� 	�  �� �  ��      F  , , 
s 6 
s � ; � ; 6 
s 6      F  , , � � � � [ � [ � � �      F  , , 
s V 
s  ;  ; V 
s V      F  , , 
s  �� 
s  � ;  � ;  �� 
s  ��      F  , , �  �f �  �. 	�  �. 	�  �f �  �f      F  , ,   ��   � �  � �  ��   ��      F  , , �  �f �  �. [  �. [  �f �  �f      F  , ,  �  n � n � �  �      F  , , 
s  � 
s  �� ;  �� ;  � 
s  �      F  , ,      � �  � �           F  , , �  � �  �^ [  �^ [  � �  �      F  , , � � � � [ � [ � � �      F  , , �  �� �  �N [  �N [  �� �  ��      F  , , 
s  �v 
s  �> ;  �> ;  �v 
s  �v      F  , , �  � �  �� [  �� [  � �  �      F  , ,   �   �^ �  �^ �  �   �      F  , , �   �  � 	�  � 	�   �        F  , , 
s  �F 
s  � ;  � ;  �F 
s  �F      F  , , � � � n [ n [ � � �      F  , , 
s  �� 
s  �N ;  �N ;  �� 
s  ��      F  , , � V �  	�  	� V � V      F  , , 
s  �� 
s  �� ;  �� ;  �� 
s  ��      F  , , 
s  �f 
s  �. ;  �. ;  �f 
s  �f      F  , , �  � �  �� 	�  �� 	�  � �  �      F  , , �  �� �  �~ 	�  �~ 	�  �� �  ��      F  , , 
s  � 
s  �^ ;  �^ ;  � 
s  �      F  , , �   �  � [  � [   �        F  , ,   �&   �� �  �� �  �&   �&      F  , , 
s  �� 
s  �� ;  �� ;  �� 
s  ��      F  , ,   �   �� �  �� �  �   �      F  , , �  �� �  �� [  �� [  �� �  ��      F  , , �  �� �  � 	�  � 	�  �� �  ��      F  , ,   ��   �N �  �N �  ��   ��      F  , , �  �F �  � [  � [  �F �  �F      F  , , �  �� �  �~ [  �~ [  �� �  ��      F  , , �  �& �  �� [  �� [  �& �  �&      F  , , 
s � 
s � ; � ; � 
s �      F  , , � � � n 	� n 	� � � �      F  , ,   ��   �~ �  �~ �  ��   ��      F  , ,   �F   � �  � �  �F   �F      F  , ,   ��   �� �  �� �  ��   ��      F  , , �  �& �  �� 	�  �� 	�  �& �  �&      F  , , � � � � 	� � 	� � � �      F  , ,   �v   �> �  �> �  �v   �v      F  , , � 6 � � [ � [ 6 � 6      F  , , �  �v �  �> [  �> [  �v �  �v      F  , , � V �  [  [ V � V      F  , , 
s   
s  � ;  � ;   
s        F  , ,  V   �  � V  V      F  , , �  �� �  �� [  �� [  �� �  ��      F  , ,  �  � � � � �  �      F  , , 
s  �& 
s  �� ;  �� ;  �& 
s  �&      F  , ,  6  � � � � 6  6      F  , , 
s � 
s n ; n ; � 
s �      F  , , �  �� �  �N 	�  �N 	�  �� �  ��      F  , , �  �F �  � 	�  � 	�  �F �  �F      E  , , �7 K� �7 La �� La �� K� �7 K�      E  , , �7 J	 �7 J� �� J� �� J	 �7 J	      E  , , �< Y2 �< Y� � Y� � Y2 �< Y2      E  , , �< W� �< Xj � Xj � W� �< W�      E  , , 
s 3� 
s 4� ; 4� ; 3� 
s 3�      E  , ,  3�  4� � 4� � 3�  3�      E  , , � 3� � 4� [ 4� [ 3� � 3�      E  , , � 3� � 4� 	� 4� 	� 3� � 3�      E  , , � �& � �� [ �� [ �& � �&      E  , , 
s �& 
s �� ; �� ; �& 
s �&      E  , ,  �&  �� � �� � �&  �&      E  , , � �& � �� 	� �� 	� �& � �&      E  , , � �f � �. [ �. [ �f � �f      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , , � �� � �� [ �� [ �� � ��      E  , , 
s �6 
s �� ; �� ; �6 
s �6      E  , , � �F � � [ � [ �F � �F      E  , , 
s �� 
s �n ; �n ; �� 
s ��      E  , , � �� � �~ [ �~ [ �� � ��      E  , , 
s � 
s �� ; �� ; � 
s �      E  , , � �� � �N [ �N [ �� � ��      E  , , 
s �� 
s �N ; �N ; �� 
s ��      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , , 
s �f 
s �. ; �. ; �f 
s �f      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , , 
s �F 
s � ; � ; �F 
s �F      E  , , 
s �� 
s �~ ; �~ ; �� 
s ��      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , ,  ��  �~ � �~ � ��  ��      E  , ,  �&  �� � �� � �&  �&      E  , ,  ��  �^ � �^ � ��  ��      E  , ,  �  �� � �� � �  �      E  , ,  �v  �> � �> � �v  �v      E  , ,  ��  �� � �� � ��  ��      E  , ,  �V  � � � � �V  �V      E  , , � �� � �~ 	� �~ 	� �� � ��      E  , ,  ��  �� � �� � ��  ��      E  , , � �& � �� 	� �� 	� �& � �&      E  , ,  �6  �� � �� � �6  �6      E  , , � �� � �^ 	� �^ 	� �� � ��      E  , ,  ��  �n � �n � ��  ��      E  , , � � � �� 	� �� 	� � � �      E  , ,  �  �� � �� � �  �      E  , , � �v � �> 	� �> 	� �v � �v      E  , ,  ��  �N � �N � ��  ��      E  , , � �� � �� 	� �� 	� �� � ��      E  , ,  ��  �� � �� � ��  ��      E  , , � �V � � 	� � 	� �V � �V      E  , , 
s �v 
s �> ; �> ; �v 
s �v      E  , ,  �f  �. � �. � �f  �f      E  , , � �� � �� 	� �� 	� �� � ��      E  , ,  ��  �� � �� � ��  ��      E  , , � �6 � �� 	� �� 	� �6 � �6      E  , ,  �F  � � � � �F  �F      E  , , � �� � �n 	� �n 	� �� � ��      E  , ,  ��  �~ � �~ � ��  ��      E  , , � � � �� 	� �� 	� � � �      E  , , � �� � �� [ �� [ �� � ��      E  , , � �� � �N 	� �N 	� �� � ��      E  , , � �� � �� 	� �� 	� �� � ��      E  , , � �f � �. 	� �. 	� �f � �f      E  , , � �� � �� 	� �� 	� �� � ��      E  , , � �F � � 	� � 	� �F � �F      E  , , � �� � �~ [ �~ [ �� � ��      E  , , � �� � �~ 	� �~ 	� �� � ��      E  , , � �& � �� [ �� [ �& � �&      E  , , 
s �V 
s � ; � ; �V 
s �V      E  , , � �� � �^ [ �^ [ �� � ��      E  , , � � � �� [ �� [ � � �      E  , , � �v � �> [ �> [ �v � �v      E  , , � �� � �� [ �� [ �� � ��      E  , , � �V � � [ � [ �V � �V      E  , , 
s �� 
s �~ ; �~ ; �� 
s ��      E  , , � �� � �� [ �� [ �� � ��      E  , , 
s �& 
s �� ; �� ; �& 
s �&      E  , , � �6 � �� [ �� [ �6 � �6      E  , , 
s �� 
s �^ ; �^ ; �� 
s ��      E  , , � �� � �n [ �n [ �� � ��      E  , , 
s � 
s �� ; �� ; � 
s �      E  , , � � � �� [ �� [ � � �      E  , , 
s oF 
s p ; p ; oF 
s oF      E  , , � p� � q� 	� q� 	� p� � p�      E  , , � {� � |� [ |� [ {� � {�      E  , , 
s m� 
s n~ ; n~ ; m� 
s m�      E  , , � z6 � z� [ z� [ z6 � z6      E  , , � u� � vN 	� vN 	� u� � u�      E  , , 
s l& 
s l� ; l� ; l& 
s l&      E  , , � w � w� 	� w� 	� w � w      E  , , � x� � yn [ yn [ x� � x�      E  , , 
s j� 
s k^ ; k^ ; j� 
s j�      E  , , 
s �� 
s �^ ; �^ ; �� 
s ��      E  , , � w � w� [ w� [ w � w      E  , , 
s � 
s �� ; �� ; � 
s �      E  , , � u� � vN [ vN [ u� � u�      E  , , 
s �v 
s �> ; �> ; �v 
s �v      E  , , � s� � t� [ t� [ s� � s�      E  , , � rf � s. [ s. [ rf � rf      E  , , 
s ~� 
s � ; � ; ~� 
s ~�      E  , , � p� � q� [ q� [ p� � p�      E  , , 
s }V 
s ~ ; ~ ; }V 
s }V      E  , , � l& � l� 	� l� 	� l& � l&      E  , , � oF � p [ p [ oF � oF      E  , , 
s {� 
s |� ; |� ; {� 
s {�      E  , ,  ��  �^ � �^ � ��  ��      E  , , � rf � s. 	� s. 	� rf � rf      E  , ,  �  �� � �� � �  �      E  , , � m� � n~ [ n~ [ m� � m�      E  , ,  �v  �> � �> � �v  �v      E  , , 
s z6 
s z� ; z� ; z6 
s z6      E  , ,  ~�  � � � � ~�  ~�      E  , , � l& � l� [ l� [ l& � l&      E  , ,  }V  ~ � ~ � }V  }V      E  , , � �� � �^ [ �^ [ �� � ��      E  , , � j� � k^ [ k^ [ j� � j�      E  , ,  {�  |� � |� � {�  {�      E  , , 
s x� 
s yn ; yn ; x� 
s x�      E  , , � j� � k^ 	� k^ 	� j� � j�      E  , ,  z6  z� � z� � z6  z6      E  , , 
s w 
s w� ; w� ; w 
s w      E  , ,  l&  l� � l� � l&  l&      E  , , � �� � �^ 	� �^ 	� �� � ��      E  , ,  x�  yn � yn � x�  x�      E  , , � oF � p 	� p 	� oF � oF      E  , , � � � �� 	� �� 	� � � �      E  , ,  w  w� � w� � w  w      E  , , 
s u� 
s vN ; vN ; u� 
s u�      E  , , � �v � �> 	� �> 	� �v � �v      E  , ,  u�  vN � vN � u�  u�      E  , , � � � �� [ �� [ � � �      E  , , � ~� � � 	� � 	� ~� � ~�      E  , ,  s�  t� � t� � s�  s�      E  , , 
s s� 
s t� ; t� ; s� 
s s�      E  , , � }V � ~ 	� ~ 	� }V � }V      E  , , � s� � t� 	� t� 	� s� � s�      E  , ,  rf  s. � s. � rf  rf      E  , , � �v � �> [ �> [ �v � �v      E  , , � {� � |� 	� |� 	� {� � {�      E  , , 
s rf 
s s. ; s. ; rf 
s rf      E  , ,  p�  q� � q� � p�  p�      E  , ,  j�  k^ � k^ � j�  j�      E  , , � z6 � z� 	� z� 	� z6 � z6      E  , , � ~� � � [ � [ ~� � ~�      E  , ,  oF  p � p � oF  oF      E  , , 
s p� 
s q� ; q� ; p� 
s p�      E  , , � x� � yn 	� yn 	� x� � x�      E  , , � m� � n~ 	� n~ 	� m� � m�      E  , ,  m�  n~ � n~ � m�  m�      E  , , � }V � ~ [ ~ [ }V � }V      E  , ,  Nv  O> � O> � Nv  Nv      E  , , � Nv � O> [ O> [ Nv � Nv      E  , , 
s Nv 
s O> ; O> ; Nv 
s Nv      E  , , � Nv � O> 	� O> 	� Nv � Nv      E  , , � ^ � ^� [ ^� [ ^ � ^      E  , , � a6 � a� 	� a� 	� a6 � a6      E  , ,  dV  e � e � dV  dV      E  , , � _� � `n [ `n [ _� � _�      E  , , � b� � c� [ c� [ b� � b�      E  , , � _� � `n 	� `n 	� _� � _�      E  , ,  VF  W � W � VF  VF      E  , , � a6 � a� [ a� [ a6 � a6      E  , ,  S&  S� � S� � S&  S&      E  , , � \� � ]N [ ]N [ \� � \�      E  , , � i � i� 	� i� 	� i � i      E  , , � Z� � [� [ [� [ Z� � Z�      E  , , � ^ � ^� 	� ^� 	� ^ � ^      E  , ,  Q�  R^ � R^ � Q�  Q�      E  , , � Yf � Z. [ Z. [ Yf � Yf      E  , ,  P  P� � P� � P  P      E  , , � \� � ]N 	� ]N 	� \� � \�      E  , , � W� � X� [ X� [ W� � W�      E  , ,  ^  ^� � ^� � ^  ^      E  , , 
s i 
s i� ; i� ; i 
s i      E  , ,  T�  U~ � U~ � T�  T�      E  , , � VF � W [ W [ VF � VF      E  , , � gv � h> 	� h> 	� gv � gv      E  , , 
s gv 
s h> ; h> ; gv 
s gv      E  , , � T� � U~ [ U~ [ T� � T�      E  , , � Z� � [� 	� [� 	� Z� � Z�      E  , , � S& � S� [ S� [ S& � S&      E  , , 
s e� 
s f� ; f� ; e� 
s e�      E  , , � Q� � R^ [ R^ [ Q� � Q�      E  , , 
s dV 
s e ; e ; dV 
s dV      E  , ,  \�  ]N � ]N � \�  \�      E  , , � P � P� [ P� [ P � P      E  , , � Yf � Z. 	� Z. 	� Yf � Yf      E  , , 
s b� 
s c� ; c� ; b� 
s b�      E  , ,  b�  c� � c� � b�  b�      E  , ,  _�  `n � `n � _�  _�      E  , , 
s a6 
s a� ; a� ; a6 
s a6      E  , , � e� � f� 	� f� 	� e� � e�      E  , , 
s _� 
s `n ; `n ; _� 
s _�      E  , , � W� � X� 	� X� 	� W� � W�      E  , , 
s ^ 
s ^� ; ^� ; ^ 
s ^      E  , ,  e�  f� � f� � e�  e�      E  , ,  Z�  [� � [� � Z�  Z�      E  , , 
s \� 
s ]N ; ]N ; \� 
s \�      E  , ,  i  i� � i� � i  i      E  , , 
s Z� 
s [� ; [� ; Z� 
s Z�      E  , , � VF � W 	� W 	� VF � VF      E  , , � dV � e 	� e 	� dV � dV      E  , , 
s Yf 
s Z. ; Z. ; Yf 
s Yf      E  , ,  Yf  Z. � Z. � Yf  Yf      E  , , � i � i� [ i� [ i � i      E  , , 
s W� 
s X� ; X� ; W� 
s W�      E  , , � T� � U~ 	� U~ 	� T� � T�      E  , ,  gv  h> � h> � gv  gv      E  , , 
s VF 
s W ; W ; VF 
s VF      E  , , � gv � h> [ h> [ gv � gv      E  , , � S& � S� 	� S� 	� S& � S&      E  , , 
s T� 
s U~ ; U~ ; T� 
s T�      E  , ,  W�  X� � X� � W�  W�      E  , , � e� � f� [ f� [ e� � e�      E  , , 
s S& 
s S� ; S� ; S& 
s S&      E  , , � Q� � R^ 	� R^ 	� Q� � Q�      E  , , � b� � c� 	� c� 	� b� � b�      E  , , 
s Q� 
s R^ ; R^ ; Q� 
s Q�      E  , , � dV � e [ e [ dV � dV      E  , ,  a6  a� � a� � a6  a6      E  , , 
s P 
s P� ; P� ; P 
s P      E  , , � P � P� 	� P� 	� P � P      E  , , � 8� � 9^ 	� 9^ 	� 8� � 8�      E  , , 
s @f 
s A. ; A. ; @f 
s @f      E  , ,  H6  H� � H� � H6  H6      E  , , 
s =F 
s > ; > ; =F 
s =F      E  , , 
s ;� 
s <~ ; <~ ; ;� 
s ;�      E  , , � I� � J� [ J� [ I� � I�      E  , , � E � E� [ E� [ E � E      E  , , � ;� � <~ 	� <~ 	� ;� � ;�      E  , ,  7  7� � 7� � 7  7      E  , , 
s KV 
s L ; L ; KV 
s KV      E  , , 
s 7 
s 7� ; 7� ; 7 
s 7      E  , ,  =F  > � > � =F  =F      E  , , � 7 � 7� 	� 7� 	� 7 � 7      E  , , � =F � > [ > [ =F � =F      E  , , � C� � DN [ DN [ C� � C�      E  , ,  I�  J� � J� � I�  I�      E  , , � C� � DN 	� DN 	� C� � C�      E  , , � 7 � 7� [ 7� [ 7 � 7      E  , , 
s :& 
s :� ; :� ; :& 
s :&      E  , ,  F�  Gn � Gn � F�  F�      E  , , � A� � B� [ B� [ A� � A�      E  , , � 5v � 6> 	� 6> 	� 5v � 5v      E  , , 
s H6 
s H� ; H� ; H6 
s H6      E  , , 
s E 
s E� ; E� ; E 
s E      E  , , � H6 � H� 	� H� 	� H6 � H6      E  , , 
s >� 
s ?� ; ?� ; >� 
s >�      E  , , � @f � A. [ A. [ @f � @f      E  , , � A� � B� 	� B� 	� A� � A�      E  , ,  E  E� � E� � E  E      E  , ,  L�  M� � M� � L�  L�      E  , , 
s C� 
s DN ; DN ; C� 
s C�      E  , , � ;� � <~ [ <~ [ ;� � ;�      E  , , 
s 5v 
s 6> ; 6> ; 5v 
s 5v      E  , , � L� � M� 	� M� 	� L� � L�      E  , ,  C�  DN � DN � C�  C�      E  , , � @f � A. 	� A. 	� @f � @f      E  , ,  5v  6> � 6> � 5v  5v      E  , , � 5v � 6> [ 6> [ 5v � 5v      E  , ,  ;�  <~ � <~ � ;�  ;�      E  , ,  A�  B� � B� � A�  A�      E  , , � E � E� 	� E� 	� E � E      E  , , � F� � Gn 	� Gn 	� F� � F�      E  , ,  >�  ?� � ?� � >�  >�      E  , , � >� � ?� 	� ?� 	� >� � >�      E  , ,  :&  :� � :� � :&  :&      E  , ,  KV  L � L � KV  KV      E  , , � >� � ?� [ ?� [ >� � >�      E  , ,  8�  9^ � 9^ � 8�  8�      E  , , � :& � :� [ :� [ :& � :&      E  , ,  @f  A. � A. � @f  @f      E  , , 
s I� 
s J� ; J� ; I� 
s I�      E  , , � L� � M� [ M� [ L� � L�      E  , , � F� � Gn [ Gn [ F� � F�      E  , , � 8� � 9^ [ 9^ [ 8� � 8�      E  , , 
s L� 
s M� ; M� ; L� 
s L�      E  , , � =F � > 	� > 	� =F � =F      E  , , � I� � J� 	� J� 	� I� � I�      E  , , 
s A� 
s B� ; B� ; A� 
s A�      E  , , � KV � L 	� L 	� KV � KV      E  , , 
s F� 
s Gn ; Gn ; F� 
s F�      E  , , � H6 � H� [ H� [ H6 � H6      E  , , � KV � L [ L [ KV � KV      E  , , � :& � :� 	� :� 	� :& � :&      E  , , 
s 8� 
s 9^ ; 9^ ; 8� 
s 8�      E  , , L |� L }] L� }] L� |� L |�      E  , , M� |� M� }] N� }] N� |� M� |�      E  , , O� |� O� }] PR }] PR |� O� |�      E  , , QL |� QL }] R }] R |� QL |�      E  , , S |� S }] S� }] S� |� S |�      E  , , � �� � �p J �p J �� � ��      E  , ,  ��  �p � �p � ��  ��      E  , , � �� � �p j �p j �� � ��      E  , , 2 �� 2 �p � �p � �� 2 ��      E  , , � �� � �p � �p � �� � ��      E  , , R �� R �p  �p  �� R ��      E  , , � �� � �p � �p � �� � ��      E  , , r �� r �p : �p : �� r ��      E  , ,  ��  �p � �p � ��  ��      E  , , � �� � �p Z �p Z �� � ��      E  , , " �� " �p � �p � �� " ��      E  , , � �� � �p z �p z �� � ��      E  , ,  B ��  B �p !
 �p !
 ��  B ��      E  , , !� �� !� �p "� �p "� �� !� ��      E  , , #b �� #b �p $* �p $* �� #b ��      E  , , $� �� $� �p %� �p %� �� $� ��      E  , , &� �� &� �p 'J �p 'J �� &� ��      E  , , ( �� ( �p (� �p (� �� ( ��      E  , , )� �� )� �p *j �p *j �� )� ��      E  , , +2 �� +2 �p +� �p +� �� +2 ��      E  , , ,� �� ,� �p -� �p -� �� ,� ��      E  , , .R �� .R �p / �p / �� .R ��      E  , , /� �� /� �p 0� �p 0� �� /� ��      E  , , 1r �� 1r �p 2: �p 2: �� 1r ��      E  , , 3 �� 3 �p 3� �p 3� �� 3 ��      E  , , 4� �� 4� �p 5Z �p 5Z �� 4� ��      E  , , 6" �� 6" �p 6� �p 6� �� 6" ��      E  , , 7� �� 7� �p 8z �p 8z �� 7� ��      E  , , � �� � �p z �p z �� � ��      E  , , B �� B �p 
 �p 
 �� B ��      E  , , � �� � �p 	� �p 	� �� � ��      E  , , 
b �� 
b �p * �p * �� 
b ��      E  , , � �� � �p � �p � �� � ��      E  , , �� �� �� �p �j �p �j �� �� ��      E  , , �2 �� �2 �p �� �p �� �� �2 ��      E  , , �� �� �� �p �� �p �� �� �� ��      E  , , �R �� �R �p � �p � �� �R ��      E  , , �� �� �� �p �� �p �� �� �� ��      E  , , �r �� �r �p  : �p  : �� �r ��      E  , ,  ��  �p � �p � ��  ��      E  , , � �� � �p Z �p Z �� � ��      E  , , " �� " �p � �p � �� " ��      E  , , .� ?9 .� @ /� @ /� ?9 .� ?9      E  , , -V ?9 -V @ . @ . ?9 -V ?9      E  , , .� @� .� A� /� A� /� @� .� @�      E  , , -V @� -V A� . A� . @� -V @�      E  , , .� BY .� C! /� C! /� BY .� BY      E  , , -V BY -V C! . C! . BY -V BY      E  , , .� C� .� D� /� D� /� C� .� C�      E  , , -V C� -V D� . D� . C� -V C�      E  , , .� Ey .� FA /� FA /� Ey .� Ey      E  , , -V Ey -V FA . FA . Ey -V Ey      E  , , .� G	 .� G� /� G� /� G	 .� G	      E  , , -V G	 -V G� . G� . G	 -V G	      E  , , .� H� .� Ia /� Ia /� H� .� H�      E  , , -V H� -V Ia . Ia . H� -V H�      E  , , w J	 w J� ? J� ? J	 w J	      E  , , � K� � La � La � K� � K�      E  , , � J	 � J� � J� � J	 � J	      E  , , W K� W La  La  K� W K�      E  , , W J	 W J�  J�  J	 W J	      E  , , � K� � La � La � K� � K�      E  , , � J	 � J� � J� � J	 � J	      E  , , 7 K� 7 La � La � K� 7 K�      E  , , 7 J	 7 J� � J� � J	 7 J	      E  , , 	� K� 	� La 
o La 
o K� 	� K�      E  , , 	� J	 	� J� 
o J� 
o J	 	� J	      E  , ,  K�  La � La � K�  K�      E  , ,  J	  J� � J� � J	  J	      E  , , � K� � La O La O K� � K�      E  , , � J	 � J� O J� O J	 � J	      E  , , � K� � La � La � K� � K�      E  , , � J	 � J� � J� � J	 � J	      E  , , g K� g La / La / K� g K�      E  , , g J	 g J� / J� / J	 g J	      E  , , � K� � La � La � K� � K�      E  , , � J	 � J� � J� � J	 � J	      E  , ,  G K�  G La  La  K�  G K�      E  , ,  G J	  G J�  J�  J	  G J	      E  , , �� K� �� La � La � K� �� K�      E  , , �� J	 �� J� � J� � J	 �� J	      E  , , �' K� �' La �� La �� K� �' K�      E  , , �' J	 �' J� �� J� �� J	 �' J	      E  , , �� K� �� La �_ La �_ K� �� K�      E  , , �� J	 �� J� �_ J� �_ J	 �� J	      E  , , � K� � La �� La �� K� � K�      E  , , � J	 � J� �� J� �� J	 � J	      E  , , �w K� �w La �? La �? K� �w K�      E  , , �w J	 �w J� �? J� �? J	 �w J	      E  , , �� K� �� La �� La �� K� �� K�      E  , , �� J	 �� J� �� J� �� J	 �� J	      E  , , �W K� �W La � La � K� �W K�      E  , , �W J	 �W J� � J� � J	 �W J	      E  , , �� K� �� La � La � K� �� K�      E  , , �� J	 �� J� � J� � J	 �� J	      E  , , .� 4I .� 5 /� 5 /� 4I .� 4I      E  , , -V 4I -V 5 . 5 . 4I -V 4I      E  , , ! K� ! La !� La !� K� ! K�      E  , , ! J	 ! J� !� J� !� J	 ! J	      E  , , � K� � La  O La  O K� � K�      E  , , � J	 � J�  O J�  O J	 � J	      E  , , � K� � La � La � K� � K�      E  , , � J	 � J� � J� � J	 � J	      E  , , g K� g La / La / K� g K�      E  , , g J	 g J� / J� / J	 g J	      E  , , � K� � La � La � K� � K�      E  , , � J	 � J� � J� � J	 � J	      E  , , G K� G La  La  K� G K�      E  , , G J	 G J�  J�  J	 G J	      E  , , � K� � La  La  K� � K�      E  , , � J	 � J�  J�  J	 � J	      E  , , ' K� ' La � La � K� ' K�      E  , , ' J	 ' J� � J� � J	 ' J	      E  , , � K� � La _ La _ K� � K�      E  , , � J	 � J� _ J� _ J	 � J	      E  , ,  K�  La � La � K�  K�      E  , ,  J	  J� � J� � J	  J	      E  , , w K� w La ? La ? K� w K�      E  , , .� 5� .� 6� /� 6� /� 5� .� 5�      E  , , -V 5� -V 6� . 6� . 5� -V 5�      E  , , .� 7i .� 81 /� 81 /� 7i .� 7i      E  , , -V 7i -V 81 . 81 . 7i -V 7i      E  , , .� 8� .� 9� /� 9� /� 8� .� 8�      E  , , -V 8� -V 9� . 9� . 8� -V 8�      E  , , .� :� .� ;Q /� ;Q /� :� .� :�      E  , , -V :� -V ;Q . ;Q . :� -V :�      E  , , .� < .� <� /� <� /� < .� <      E  , , -V < -V <� . <� . < -V <      E  , , .� =� .� >q /� >q /� =� .� =�      E  , , -V =� -V >q . >q . =� -V =�      E  , , .� �� .� �a /� �a /� �� .� ��      E  , , -V �� -V �a . �a . �� -V ��      E  , , .� Y .� ! /� ! /� Y .� Y      E  , , -V Y -V ! . ! . Y -V Y      E  , , .� � .� � /� � /� � .� �      E  , , -V � -V � . � . � -V �      E  , , .� y .� A /� A /� y .� y      E  , , -V y -V A . A . y -V y      E  , , .� 	 .� � /� � /� 	 .� 	      E  , , -V 	 -V � . � . 	 -V 	      E  , , .� � .� a /� a /� � .� �      E  , , -V � -V a . a . � -V �      E  , , .� ) .� � /� � /� ) .� )      E  , , -V ) -V � . � . ) -V )      E  , , .� � .� � /� � /� � .� �      E  , , -V � -V � . � . � -V �      E  , , .� I .�  /�  /� I .� I      E  , , -V I -V  .  . I -V I      E  , , .� � .� � /� � /� � .� �      E  , , -V � -V � . � . � -V �      E  , , .� i .� 1 /� 1 /� i .� i      E  , , -V i -V 1 . 1 . i -V i      E  , , .� � .�  � /�  � /� � .� �      E  , , -V � -V  � .  � . � -V �      E  , , .� !� .� "Q /� "Q /� !� .� !�      E  , , -V !� -V "Q . "Q . !� -V !�      E  , , .� # .� #� /� #� /� # .� #      E  , , -V # -V #� . #� . # -V #      E  , , .� $� .� %q /� %q /� $� .� $�      E  , , -V $� -V %q . %q . $� -V $�      E  , , .� &9 .� ' /� ' /� &9 .� &9      E  , , -V &9 -V ' . ' . &9 -V &9      E  , , .� '� .� (� /� (� /� '� .� '�      E  , , -V '� -V (� . (� . '� -V '�      E  , , .� )Y .� *! /� *! /� )Y .� )Y      E  , , -V )Y -V *! . *! . )Y -V )Y      E  , , .� *� .� +� /� +� /� *� .� *�      E  , , -V *� -V +� . +� . *� -V *�      E  , , .� ,y .� -A /� -A /� ,y .� ,y      E  , , -V ,y -V -A . -A . ,y -V ,y      E  , , .� .	 .� .� /� .� /� .	 .� .	      E  , , -V .	 -V .� . .� . .	 -V .	      E  , , .� /� .� 0a /� 0a /� /� .� /�      E  , , -V /� -V 0a . 0a . /� -V /�      E  , , .� 1) .� 1� /� 1� /� 1) .� 1)      E  , , -V 1) -V 1� . 1� . 1) -V 1)      E  , , .� 2� .� 3� /� 3� /� 2� .� 2�      E  , , -V 2� -V 3� . 3� . 2� -V 2�      E  , , .� � .� � /� � /� � .� �      E  , , -V � -V � . � . � -V �      E  , , .� �) .� �� /� �� /� �) .� �)      E  , , -V �) -V �� . �� . �) -V �)      E  , , .�  � .� � /� � /�  � .�  �      E  , , -V  � -V � . � .  � -V  �      E  , , .� I .�  /�  /� I .� I      E  , , -V I -V  .  . I -V I      E  , , .� � .� � /� � /� � .� �      E  , , -V � -V � . � . � -V �      E  , , .� i .� 1 /� 1 /� i .� i      E  , , -V i -V 1 . 1 . i -V i      E  , , .� � .� � /� � /� � .� �      E  , , -V � -V � . � . � -V �      E  , , .� � .� 	Q /� 	Q /� � .� �      E  , , -V � -V 	Q . 	Q . � -V �      E  , , .� 
 .� 
� /� 
� /� 
 .� 
      E  , , -V 
 -V 
� . 
� . 
 -V 
      E  , , .� � .� q /� q /� � .� �      E  , , -V � -V q . q . � -V �      E  , , .� 9 .�  /�  /� 9 .� 9      E  , , -V 9 -V  .  . 9 -V 9      E  , , -V �� -V � . � . �� -V ��      E  , , .� �y .� �A /� �A /� �y .� �y      E  , , -V �y -V �A . �A . �y -V �y      E  , , .� �	 .� �� /� �� /� �	 .� �	      E  , , -V �	 -V �� . �� . �	 -V �	      E  , , .� � .� �a /� �a /� � .� �      E  , , -V � -V �a . �a . � -V �      E  , , .� �) .� �� /� �� /� �) .� �)      E  , , -V �) -V �� . �� . �) -V �)      E  , , .� � .� � /� � /� � .� �      E  , , -V � -V � . � . � -V �      E  , , .� �I .� � /� � /� �I .� �I      E  , , -V �I -V � . � . �I -V �I      E  , , .� �� .� � /� � /� �� .� ��      E  , , -V �� -V � . � . �� -V ��      E  , , .� �i .� �1 /� �1 /� �i .� �i      E  , , -V �i -V �1 . �1 . �i -V �i      E  , , .� �� .� �� /� �� /� �� .� ��      E  , , .� �y .� �A /� �A /� �y .� �y      E  , , -V �y -V �A . �A . �y -V �y      E  , , .� �	 .� �� /� �� /� �	 .� �	      E  , , -V �	 -V �� . �� . �	 -V �	      E  , , .� ˙ .� �a /� �a /� ˙ .� ˙      E  , , -V ˙ -V �a . �a . ˙ -V ˙      E  , , .� �) .� �� /� �� /� �) .� �)      E  , , -V �) -V �� . �� . �) -V �)      E  , , .� ι .� ρ /� ρ /� ι .� ι      E  , , -V ι -V ρ . ρ . ι -V ι      E  , , .� �I .� � /� � /� �I .� �I      E  , , -V �I -V � . � . �I -V �I      E  , , .� �� .� ҡ /� ҡ /� �� .� ��      E  , , -V �� -V ҡ . ҡ . �� -V ��      E  , , .� �i .� �1 /� �1 /� �i .� �i      E  , , -V �i -V �1 . �1 . �i -V �i      E  , , .� �� .� �� /� �� /� �� .� ��      E  , , -V �� -V �� . �� . �� -V ��      E  , , .� ։ .� �Q /� �Q /� ։ .� ։      E  , , -V ։ -V �Q . �Q . ։ -V ։      E  , , .� � .� �� /� �� /� � .� �      E  , , -V � -V �� . �� . � -V �      E  , , .� ٩ .� �q /� �q /� ٩ .� ٩      E  , , -V ٩ -V �q . �q . ٩ -V ٩      E  , , .� �9 .� � /� � /� �9 .� �9      E  , , -V �9 -V � . � . �9 -V �9      E  , , .� �	 .� �� /� �� /� �	 .� �	      E  , , -V �	 -V �� . �� . �	 -V �	      E  , , .� �� .� ݑ /� ݑ /� �� .� ��      E  , , -V �� -V ݑ . ݑ . �� -V ��      E  , , .� �Y .� �! /� �! /� �Y .� �Y      E  , , -V �Y -V �! . �! . �Y -V �Y      E  , , .� �� .� � /� � /� �� .� ��      E  , , .� � .� �q /� �q /� � .� �      E  , , -V � -V �q . �q . � -V �      E  , , .� �9 .� � /� � /� �9 .� �9      E  , , -V �9 -V � . � . �9 -V �9      E  , , .� �� .� �� /� �� /� �� .� ��      E  , , -V �� -V �� . �� . �� -V ��      E  , , .� �Y .� �! /� �! /� �Y .� �Y      E  , , -V �Y -V �! . �! . �Y -V �Y      E  , , .� �� .� �� /� �� /� �� .� ��      E  , , -V �� -V �� . �� . �� -V ��      E  , , .� �y .� �A /� �A /� �y .� �y      E  , , -V �y -V �A . �A . �y -V �y      E  , , .� � .� �Q /� �Q /� � .� �      E  , , -V � -V �Q . �Q . � -V �      E  , , .� � .� �� /� �� /� � .� �      E  , , -V � -V �� . �� . � -V �      E  , , -V �� -V �� . �� . �� -V ��      E  , , � �6 � �� 	� �� 	� �6 � �6      E  , , � �6 � �� [ �� [ �6 � �6      E  , , 
s �6 
s �� ; �� ; �6 
s �6      E  , ,  �6  �� � �� � �6  �6      E  , , 
s 0� 
s 1� ; 1� ; 0� 
s 0�      E  , ,    � � � �         E  , , �  � � [ � [  �       E  , , � V �  	�  	� V � V      E  , , � v � > [ > [ v � v      E  , , � 2V � 3 	� 3 	� 2V � 2V      E  , , � � � � [ � [ � � �      E  , , 
s � 
s � ; � ; � 
s �      E  , ,  �  � � � � �  �      E  , , � V �  [  [ V � V      E  , , � 0� � 1� 	� 1� 	� 0� � 0�      E  , , 
s /6 
s /� ; /� ; /6 
s /6      E  , , � /6 � /� 	� /� 	� /6 � /6      E  , , 
s V 
s  ;  ; V 
s V      E  , , � -� � .n 	� .n 	� -� � -�      E  , ,  V   �  � V  V      E  , , � "� � #~ 	� #~ 	� "� � "�      E  , , � 'f � (. 	� (. 	� 'f � 'f      E  , , � , � ,� 	� ,� 	� , � ,      E  , , 
s -� 
s .n ; .n ; -� 
s -�      E  , , � *� � +N 	� +N 	� *� � *�      E  , , � (� � )� 	� )� 	� (� � (�      E  , ,  �   ^ �  ^ � �  �      E  , , � � �  ^ [  ^ [ � � �      E  , , 
s v 
s > ; > ; v 
s v      E  , ,  v  > � > � v  v      E  , , �  � � 	� � 	�  �       E  , , 
s *� 
s +N ; +N ; *� 
s *�      E  , , 
s (� 
s )� ; )� ; (� 
s (�      E  , , 
s 'f 
s (. ; (. ; 'f 
s 'f      E  , , � $F � % 	� % 	� $F � $F      E  , ,  2V  3 � 3 � 2V  2V      E  , , � 2V � 3 [ 3 [ 2V � 2V      E  , ,  0�  1� � 1� � 0�  0�      E  , , � 0� � 1� [ 1� [ 0� � 0�      E  , , 
s %� 
s &� ; &� ; %� 
s %�      E  , , � v � > 	� > 	� v � v      E  , , � !& � !� 	� !� 	� !& � !&      E  , ,  /6  /� � /� � /6  /6      E  , , � /6 � /� [ /� [ /6 � /6      E  , , 
s $F 
s % ; % ; $F 
s $F      E  , ,  -�  .n � .n � -�  -�      E  , , � -� � .n [ .n [ -� � -�      E  , , � %� � &� 	� &� 	� %� � %�      E  , ,  ,  ,� � ,� � ,  ,      E  , , � , � ,� [ ,� [ , � ,      E  , , 
s "� 
s #~ ; #~ ; "� 
s "�      E  , ,  *�  +N � +N � *�  *�      E  , , � *� � +N [ +N [ *� � *�      E  , ,  (�  )� � )� � (�  (�      E  , , � (� � )� [ )� [ (� � (�      E  , , � � � � 	� � 	� � � �      E  , , 
s !& 
s !� ; !� ; !& 
s !&      E  , ,  'f  (. � (. � 'f  'f      E  , , � 'f � (. [ (. [ 'f � 'f      E  , , 
s � 
s  ^ ;  ^ ; � 
s �      E  , ,  %�  &� � &� � %�  %�      E  , , � %� � &� [ &� [ %� � %�      E  , ,  $F  % � % � $F  $F      E  , , � $F � % [ % [ $F � $F      E  , ,  "�  #~ � #~ � "�  "�      E  , , � "� � #~ [ #~ [ "� � "�      E  , , 
s  
s � ; � ;  
s       E  , , 
s 2V 
s 3 ; 3 ; 2V 
s 2V      E  , ,  !&  !� � !� � !&  !&      E  , , � !& � !� [ !� [ !& � !&      E  , , � � �  ^ 	�  ^ 	� � � �      E  , , 
s , 
s ,� ; ,� ; , 
s ,      E  , , �  V �  	�  	�  V �  V      E  , , � F �  [  [ F � F      E  , , 
s & 
s � ; � ; & 
s &      E  , ,  �  � � � � �  �      E  , ,  &  � � � � &  &      E  , , � � � � [ � [ � � �      E  , , � 6 � � 	� � 	� 6 � 6      E  , , � 	� � 
~ 	� 
~ 	� 	� � 	�      E  , , � � � n 	� n 	� � � �      E  , , � v � > [ > [ v � v      E  , , � � � � 	� � 	� � � �      E  , , 
s 6 
s � ; � ; 6 
s 6      E  , , � �� � �� [ �� [ �� � ��      E  , , �  � � [ � [  �       E  , , 
s � 
s ^ ; ^ ; � 
s �      E  , , 
s � 
s � ; � ; � 
s �      E  , , � � � � [ � [ � � �      E  , ,  �  ^ � ^ � �  �      E  , , � 6 � � [ � [ 6 � 6      E  , ,  �  � � � � �  �      E  , , �  V �  [  [  V �  V      E  , , 
s f 
s . ; . ; f 
s f      E  , , � �� � �� 	� �� 	� �� � ��      E  , , 
s v 
s > ; > ; v 
s v      E  , , � & � � [ � [ & � &      E  , , � � � n [ n [ � � �      E  , ,  f  . � . � f  f      E  , , � � � � 	� � 	� � � �      E  , , 
s  
s � ; � ;  
s       E  , , � � � N 	� N 	� � � �      E  , , �  � � [ � [  �       E  , , 
s  V 
s  ;  ;  V 
s  V      E  , , � F �  	�  	� F � F      E  , , 
s  
s � ; � ;  
s       E  , , � � � N [ N [ � � �      E  , ,   V   �  �  V   V      E  , ,    � � � �         E  , , 
s � 
s � ; � ; � 
s �      E  , , � v � > 	� > 	� v � v      E  , ,  �  � � � � �  �      E  , , � � � � [ � [ � � �      E  , , 
s � 
s N ; N ; � 
s �      E  , ,    � � � �         E  , , � � � � 	� � 	� � � �      E  , ,  �  N � N � �  �      E  , , � f � . [ . [ f � f      E  , , � � � � 	� � 	� � � �      E  , ,  v  > � > � v  v      E  , , 
s F 
s  ;  ; F 
s F      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , ,  ��  �� � �� � ��  ��      E  , , � � � ^ 	� ^ 	� � � �      E  , ,  F   �  � F  F      E  , , � � � ^ [ ^ [ � � �      E  , , �  � � 	� � 	�  �       E  , , � & � � 	� � 	� & � &      E  , ,  6  � � � � 6  6      E  , , 
s � 
s n ; n ; � 
s �      E  , , � f � . 	� . 	� f � f      E  , , � � � � [ � [ � � �      E  , , �  � � 	� � 	�  �       E  , , 
s 	� 
s 
~ ; 
~ ; 	� 
s 	�      E  , ,  	�  
~ � 
~ � 	�  	�      E  , , � 	� � 
~ [ 
~ [ 	� � 	�      E  , , 
s � 
s � ; � ; � 
s �      E  , ,  �  � � � � �  �      E  , ,  �  n � n � �  �      E  , , 
s � 
s � ; � ; � 
s �      E  , ,  �  �n � �n � �  �      E  , , � � � �n [ �n [ � � �      E  , , � � � �n 	� �n 	� � � �      E  , , 
s � 
s �n ; �n ; � 
s �      E  , , 
s � 
s �� ; �� ; � 
s �      E  , , 
s �F 
s � ; � ; �F 
s �F      E  , ,  �  �~ � �~ � �  �      E  , ,  �&  �� � �� � �&  �&      E  , , � � � �� [ �� [ � � �      E  , , � �6 � �� 	� �� 	� �6 � �6      E  , , � �f � �. 	� �. 	� �f � �f      E  , , � � � �� 	� �� 	� � � �      E  , , � �� � �� 	� �� 	� �� � ��      E  , , 
s �v 
s �> ; �> ; �v 
s �v      E  , ,  �F  � � � � �F  �F      E  , , � �& � �� 	� �� 	� �& � �&      E  , , � �F � � [ � [ �F � �F      E  , ,  �V  � � � � �V  �V      E  , ,  �v  �> � �> � �v  �v      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , , 
s �& 
s �� ; �� ; �& 
s �&      E  , , � �f � �. [ �. [ �f � �f      E  , , � �6 � �� [ �� [ �6 � �6      E  , , � �� � � 	� � 	� �� � ��      E  , , � �� � �� 	� �� 	� �� � ��      E  , ,  ��  � � � � ��  ��      E  , , � �v � �> [ �> [ �v � �v      E  , , 
s �� 
s � ; � ; �� 
s ��      E  , ,  ��  �� � �� � ��  ��      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , , � �� � �n 	� �n 	� �� � ��      E  , , � �V � � [ � [ �V � �V      E  , , � � � �~ [ �~ [ � � �      E  , , � �V � � 	� � 	� �V � �V      E  , , 
s �f 
s �. ; �. ; �f 
s �f      E  , , � � � �� 	� �� 	� � � �      E  , , 
s � 
s �� ; �� ; � 
s �      E  , , 
s �V 
s � ; � ; �V 
s �V      E  , , � �v � �> 	� �> 	� �v � �v      E  , , � �� � �� [ �� [ �� � ��      E  , , � � � �^ 	� �^ 	� � � �      E  , , 
s �6 
s �� ; �� ; �6 
s �6      E  , , 
s � 
s �^ ; �^ ; � 
s �      E  , , 
s �� 
s �n ; �n ; �� 
s ��      E  , ,  ��  �n � �n � ��  ��      E  , , � � � �� [ �� [ � � �      E  , ,  �6  �� � �� � �6  �6      E  , ,  �  �� � �� � �  �      E  , , � �� � �N 	� �N 	� �� � ��      E  , , � �F � � 	� � 	� �F � �F      E  , , 
s �� 
s �N ; �N ; �� 
s ��      E  , , � �� � � 	� � 	� �� � ��      E  , , � �� � �n [ �n [ �� � ��      E  , , � �& � �� [ �� [ �& � �&      E  , ,  ��  �N � �N � ��  ��      E  , ,  �  �� � �� � �  �      E  , , 
s �� 
s � ; � ; �� 
s ��      E  , , � � � �^ [ �^ [ � � �      E  , , � �� � �N [ �N [ �� � ��      E  , , � � � �~ 	� �~ 	� � � �      E  , , � �� � � [ � [ �� � ��      E  , ,  ��  �� � �� � ��  ��      E  , , � �� � �� [ �� [ �� � ��      E  , ,  ��  � � � � ��  ��      E  , , 
s � 
s �~ ; �~ ; � 
s �      E  , ,  �  �^ � �^ � �  �      E  , ,  �f  �. � �. � �f  �f      E  , , � �� � � [ � [ �� � ��      E  , , � �F � � 	� � 	� �F � �F      E  , , 
s � 
s �� ; �� ; � 
s �      E  , , 
s � 
s �� ; �� ; � 
s �      E  , ,  �  �� � �� � �  �      E  , , � �� � Ю [ Ю [ �� � ��      E  , , � �� � ޾ 	� ޾ 	� �� � ��      E  , , � �F � � [ � [ �F � �F      E  , , � Ԗ � �^ [ �^ [ Ԗ � Ԗ      E  , , 
s ߆ 
s �N ; �N ; ߆ 
s ߆      E  , , 
s �f 
s �. ; �. ; �f 
s �f      E  , , � �& � �� 	� �� 	� �& � �&      E  , ,  ��  ۞ � ۞ � ��  ��      E  , , 
s �F 
s � ; � ; �F 
s �F      E  , ,  �  �� � �� � �  �      E  , , � ׶ � �~ [ �~ [ ׶ � ׶      E  , ,  Ԗ  �^ � �^ � Ԗ  Ԗ      E  , , � �� � ͎ [ ͎ [ �� � ��      E  , ,  �V  � � � � �V  �V      E  , ,  ��  ޾ � ޾ � ��  ��      E  , , � � � �� [ �� [ � � �      E  , , � �v � �> [ �> [ �v � �v      E  , ,  ߆  �N � �N � ߆  ߆      E  , , 
s ɦ 
s �n ; �n ; ɦ 
s ɦ      E  , ,  ׶  �~ � �~ � ׶  ׶      E  , ,  �F  � � � � �F  �F      E  , , � �V � � 	� � 	� �V � �V      E  , , 
s �v 
s �> ; �> ; �v 
s �v      E  , , � ׶ � �~ 	� �~ 	� ׶ � ׶      E  , ,  �&  �� � �� � �&  �&      E  , ,  �  �� � �� � �  �      E  , , � ɦ � �n [ �n [ ɦ � ɦ      E  , , 
s �� 
s ޾ ; ޾ ; �� 
s ��      E  , , � �� � ͎ 	� ͎ 	� �� � ��      E  , ,  �v  �> � �> � �v  �v      E  , ,  ��  ͎ � ͎ � ��  ��      E  , , � ߆ � �N [ �N [ ߆ � ߆      E  , , � �� � Ю 	� Ю 	� �� � ��      E  , , 
s �� 
s ۞ ; ۞ ; �� 
s ��      E  , , 
s �� 
s ͎ ; ͎ ; �� 
s ��      E  , ,  �6  �� � �� � �6  �6      E  , , � �& � �� [ �� [ �& � �&      E  , , � �6 � �� 	� �� 	� �6 � �6      E  , , 
s ׶ 
s �~ ; �~ ; ׶ 
s ׶      E  , , � � � �� 	� �� 	� � � �      E  , , � �� � ۞ 	� ۞ 	� �� � ��      E  , , � �V � � [ � [ �V � �V      E  , , � �f � �. [ �. [ �f � �f      E  , , � �f � �. 	� �. 	� �f � �f      E  , , � �v � �> 	� �> 	� �v � �v      E  , , � �� � ۞ [ ۞ [ �� � ��      E  , , 
s �� 
s Ю ; Ю ; �� 
s ��      E  , , � �6 � �� [ �� [ �6 � �6      E  , , 
s �& 
s �� ; �� ; �& 
s �&      E  , , � � � �� 	� �� 	� � � �      E  , , � ɦ � �n 	� �n 	� ɦ � ɦ      E  , , 
s � 
s �� ; �� ; � 
s �      E  , , � � � �� [ �� [ � � �      E  , , 
s �6 
s �� ; �� ; �6 
s �6      E  , , � �� � ޾ [ ޾ [ �� � ��      E  , , � � � �� 	� �� 	� � � �      E  , , 
s �V 
s � ; � ; �V 
s �V      E  , , � � � �� [ �� [ � � �      E  , , � Ԗ � �^ 	� �^ 	� Ԗ � Ԗ      E  , , 
s Ԗ 
s �^ ; �^ ; Ԗ 
s Ԗ      E  , ,  ɦ  �n � �n � ɦ  ɦ      E  , ,  ��  Ю � Ю � ��  ��      E  , ,  �f  �. � �. � �f  �f      E  , , � ߆ � �N 	� �N 	� ߆ � ߆      E  , ,  �� 3�  �� 4�  � 4�  � 3�  �� 3�      E  , ,  �a 3�  �a 4�  �) 4�  �) 3�  �a 3�      E  , , �� K� �� La �� La �� K� �� K�      E  , , �� J	 �� J� �� J� �� J	 �� J	      E  , , �W K� �W La � La � K� �W K�      E  , , �W J	 �W J� � J� � J	 �W J	      E  , , �� K� �� La �� La �� K� �� K�      E  , , �� J	 �� J� �� J� �� J	 �� J	      E  , , �7 K� �7 La �� La �� K� �7 K�      E  , , �7 J	 �7 J� �� J� �� J	 �7 J	      E  , , �� K� �� La �o La �o K� �� K�      E  , , �� J	 �� J� �o J� �o J	 �� J	      E  , , � K� � La �� La �� K� � K�      E  , , � J	 � J� �� J� �� J	 � J	      E  , , �� K� �� La �O La �O K� �� K�      E  , , �� J	 �� J� �O J� �O J	 �� J	      E  , , �� K� �� La �� La �� K� �� K�      E  , , �� J	 �� J� �� J� �� J	 �� J	      E  , , �g K� �g La �/ La �/ K� �g K�      E  , , �g J	 �g J� �/ J� �/ J	 �g J	      E  , , �� K� �� La �� La �� K� �� K�      E  , , �� J	 �� J� �� J� �� J	 �� J	      E  , , �G K� �G La � La � K� �G K�      E  , , �G J	 �G J� � J� � J	 �G J	      E  , , �� K� �� La � La � K� �� K�      E  , , �� J	 �� J� � J� � J	 �� J	      E  , , �' K� �' La �� La �� K� �' K�      E  , , �' J	 �' J� �� J� �� J	 �' J	      E  , , �� K� �� La �_ La �_ K� �� K�      E  , , �� J	 �� J� �_ J� �_ J	 �� J	      E  , , � K� � La �� La �� K� � K�      E  , , � J	 � J� �� J� �� J	 � J	      E  , , �w K� �w La �? La �? K� �w K�      E  , , �w J	 �w J� �? J� �? J	 �w J	      E  , , �� K� �� La �� La �� K� �� K�      E  , , �� J	 �� J� �� J� �� J	 �� J	      E  , , �W K� �W La � La � K� �W K�      E  , , �W J	 �W J� � J� � J	 �W J	      E  , , �� K� �� La �� La �� K� �� K�      E  , , �� J	 �� J� �� J� �� J	 �� J	      E  , , �7 K� �7 La �� La �� K� �7 K�      E  , , �7 J	 �7 J� �� J� �� J	 �7 J	      E  , , �� K� �� La �o La �o K� �� K�      E  , , �� J	 �� J� �o J� �o J	 �� J	      E  , , � K� � La �� La �� K� � K�      E  , , � J	 � J� �� J� �� J	 � J	      E  , , �� K� �� La �O La �O K� �� K�      E  , , �� J	 �� J� �O J� �O J	 �� J	      E  , , �� K� �� La �� La �� K� �� K�      E  , , �� J	 �� J� �� J� �� J	 �� J	      E  , , e� Qu e� R= fU R= fU Qu e� Qu      E  , , e� S e� S� fU S� fU S e� S      E  , , g Qu g R= g� R= g� Qu g Qu      E  , , g S g S� g� S� g� S g S      E  , , h� Qu h� R= iu R= iu Qu h� Qu      E  , , h� S h� S� iu S� iu S h� S      E  , , j= Qu j= R= k R= k Qu j= Qu      E  , , j= S j= S� k S� k S j= S      E  , , k� Qu k� R= l� R= l� Qu k� Qu      E  , , k� S k� S� l� S� l� S k� S      E  , , m] Qu m] R= n% R= n% Qu m] Qu      E  , , m] S m] S� n% S� n% S m] S      E  , , n� Qu n� R= o� R= o� Qu n� Qu      E  , , n� S n� S� o� S� o� S n� S      E  , , p} Qu p} R= qE R= qE Qu p} Qu      E  , , p} S p} S� qE S� qE S p} S      E  , , � K� � La �� La �� K� � K�      E  , , � J	 � J� �� J� �� J	 � J	      E  , , �w K� �w La �? La �? K� �w K�      E  , , �w J	 �w J� �? J� �? J	 �w J	      E  , , �� K� �� La ů La ů K� �� K�      E  , , �� J	 �� J� ů J� ů J	 �� J	      E  , , �W K� �W La � La � K� �W K�      E  , , �W J	 �W J� � J� � J	 �W J	      E  , , �� K� �� La  La  K� �� K�      E  , , �� J	 �� J�  J�  J	 �� J	      E  , , �7 K� �7 La �� La �� K� �7 K�      E  , , �7 J	 �7 J� �� J� �� J	 �7 J	      E  , , �� K� �� La �o La �o K� �� K�      E  , , �� J	 �� J� �o J� �o J	 �� J	      E  , , � K� � La �� La �� K� � K�      E  , , � J	 � J� �� J� �� J	 � J	      E  , , �� K� �� La �O La �O K� �� K�      E  , , �� J	 �� J� �O J� �O J	 �� J	      E  , , �� K� �� La �� La �� K� �� K�      E  , , �� J	 �� J� �� J� �� J	 �� J	      E  , , �g K� �g La �/ La �/ K� �g K�      E  , , �g J	 �g J� �/ J� �/ J	 �g J	      E  , , �� K� �� La �� La �� K� �� K�      E  , , �� J	 �� J� �� J� �� J	 �� J	      E  , , �G K� �G La � La � K� �G K�      E  , , �G J	 �G J� � J� � J	 �G J	      E  , , �� K� �� La � La � K� �� K�      E  , , �� J	 �� J� � J� � J	 �� J	      E  , , �' K� �' La �� La �� K� �' K�      E  , , �' J	 �' J� �� J� �� J	 �' J	      E  , , �� K� �� La �_ La �_ K� �� K�      E  , , �� J	 �� J� �_ J� �_ J	 �� J	      E  , , � K� � La �� La �� K� � K�      E  , , � J	 � J� �� J� �� J	 � J	      E  , , � J	 � J� �o J� �o J	 � J	      E  , , � K� � La �� La �� K� � K�      E  , , � J	 � J� �� J� �� J	 � J	      E  , , � K� � La �O La �O K� � K�      E  , , � J	 � J� �O J� �O J	 � J	      E  , , �� K� �� La � La � K� �� K�      E  , , �� J	 �� J� � J� � J	 �� J	      E  , , �g K� �g La �/ La �/ K� �g K�      E  , , �g J	 �g J� �/ J� �/ J	 �g J	      E  , , �� K� �� La � La � K� �� K�      E  , , �� J	 �� J� � J� � J	 �� J	      E  , , �G K� �G La � La � K� �G K�      E  , , �G J	 �G J� � J� � J	 �G J	      E  , , � K� � La � La � K� � K�      E  , , � J	 � J� � J� � J	 � J	      E  , , �' K� �' La �� La �� K� �' K�      E  , , �' J	 �' J� �� J� �� J	 �' J	      E  , , � K� � La �_ La �_ K� � K�      E  , , �w K� �w La �? La �? K� �w K�      E  , , �w J	 �w J� �? J� �? J	 �w J	      E  , , �� K� �� La ӿ La ӿ K� �� K�      E  , , �� J	 �� J� ӿ J� ӿ J	 �� J	      E  , , �g K� �g La �/ La �/ K� �g K�      E  , , �g J	 �g J� �/ J� �/ J	 �g J	      E  , , �� K� �� La П La П K� �� K�      E  , , �� J	 �� J� П J� П J	 �� J	      E  , , �G K� �G La � La � K� �G K�      E  , , �G J	 �G J� � J� � J	 �G J	      E  , , ̷ K� ̷ La � La � K� ̷ K�      E  , , ̷ J	 ̷ J� � J� � J	 ̷ J	      E  , , �' K� �' La �� La �� K� �' K�      E  , , �' J	 �' J� �� J� �� J	 �' J	      E  , , ɗ K� ɗ La �_ La �_ K� ɗ K�      E  , , ɗ J	 ɗ J� �_ J� �_ J	 ɗ J	      E  , , � K� � La �o La �o K� � K�      E  , , �� K� �� La ޯ La ޯ K� �� K�      E  , , �� J	 �� J� ޯ J� ޯ J	 �� J	      E  , , �W K� �W La � La � K� �W K�      E  , , �W J	 �W J� � J� � J	 �W J	      E  , , �� K� �� La ۏ La ۏ K� �� K�      E  , , �� J	 �� J� ۏ J� ۏ J	 �� J	      E  , , �7 K� �7 La �� La �� K� �7 K�      E  , , �7 J	 �7 J� �� J� �� J	 �7 J	      E  , , ק K� ק La �o La �o K� ק K�      E  , , ק J	 ק J� �o J� �o J	 ק J	      E  , , � K� � La �� La �� K� � K�      E  , , � J	 � J� �� J� �� J	 � J	      E  , , � K� � La �� La �� K� � K�      E  , , � J	 � J� �� J� �� J	 � J	      E  , , �w K� �w La �? La �? K� �w K�      E  , , �w J	 �w J� �? J� �? J	 �w J	      E  , , � J	 � J� �_ J� �_ J	 � J	      E  , , ԇ K� ԇ La �O La �O K� ԇ K�      E  , , ԇ J	 ԇ J� �O J� �O J	 ԇ J	      E  , , � Qu � R= u R= u Qu � Qu      E  , , � S � S� u S� u S � S      E  , ,  �M Qu  �M R=  � R=  � Qu  �M Qu      E  , ,  �M S  �M S�  � S�  � S  �M S      E  , ,  �� Qu  �� R=  �� R=  �� Qu  �� Qu      E  , ,  �� S  �� S�  �� S�  �� S  �� S      E  , ,  �m Qu  �m R=  �5 R=  �5 Qu  �m Qu      E  , ,  �m S  �m S�  �5 S�  �5 S  �m S      E  , ,  �� Qu  �� R=  � R=  � Qu  �� Qu      E  , ,  �� S  �� S�  � S�  � S  �� S      E  , , � Qu � R= U R= U Qu � Qu      E  , , � S � S� U S� U S � S      E  , ,  Qu  R= � R= � Qu  Qu      E  , ,  S  S� � S� � S  S      E  , , � Qu � R= u R= u Qu � Qu      E  , , � S � S� u S� u S � S      E  , , = Qu = R=  R=  Qu = Qu      E  , , = S = S�  S�  S = S      E  , , � Qu � R= � R= � Qu � Qu      E  , , � S � S� � S� � S � S      E  , , 	] Qu 	] R= 
% R= 
% Qu 	] Qu      E  , , 	] S 	] S� 
% S� 
% S 	] S      E  , , 
� Qu 
� R= � R= � Qu 
� Qu      E  , , 
� S 
� S� � S� � S 
� S      E  , , } Qu } R= E R= E Qu } Qu      E  , , } S } S� E S� E S } S      E  , ,  Qu  R= � R= � Qu  Qu      E  , ,  S  S� � S� � S  S      E  , , � Qu � R= e R= e Qu � Qu      E  , , � S � S� e S� e S � S      E  , , - Qu - R= � R= � Qu - Qu      E  , , - S - S� � S� � S - S      E  , , � Qu � R= � R= � Qu � Qu      E  , , � S � S� � S� � S � S      E  , , M Qu M R=  R=  Qu M Qu      E  , , M S M S�  S�  S M S      E  , , � Qu � R= � R= � Qu � Qu      E  , , m Qu m R= 5 R= 5 Qu m Qu      E  , , m S m S� 5 S� 5 S m S      E  , , � Qu � R= � R= � Qu � Qu      E  , , � S � S� � S� � S � S      E  , , � Qu � R= U R= U Qu � Qu      E  , , � S � S� U S� U S � S      E  , ,  Qu  R= � R= � Qu  Qu      E  , ,  S  S� � S� � S  S      E  , , � S � S� � S� � S � S      E  , ,  �� Qu  �� R=  �� R=  �� Qu  �� Qu      E  , ,  �� S  �� S�  �� S�  �� S  �� S      E  , ,  �] Qu  �] R=  �% R=  �% Qu  �] Qu      E  , ,  �] S  �] S�  �% S�  �% S  �] S      E  , ,  �� Qu  �� R=  ٵ R=  ٵ Qu  �� Qu      E  , ,  �� S  �� S�  ٵ S�  ٵ S  �� S      E  , ,  �} Qu  �} R=  �E R=  �E Qu  �} Qu      E  , ,  �} S  �} S�  �E S�  �E S  �} S      E  , ,  � Qu  � R=  �� R=  �� Qu  � Qu      E  , ,  � S  � S�  �� S�  �� S  � S      E  , ,  ݝ Qu  ݝ R=  �e R=  �e Qu  ݝ Qu      E  , ,  ݝ S  ݝ S�  �e S�  �e S  ݝ S      E  , ,  �- Qu  �- R=  �� R=  �� Qu  �- Qu      E  , ,  �- S  �- S�  �� S�  �� S  �- S      E  , ,  � Qu  � R=  � R=  � Qu  � Qu      E  , ,  � S  � S�  � S�  � S  � S      E  , ,  �M Qu  �M R=  � R=  � Qu  �M Qu      E  , ,  �M S  �M S�  � S�  � S  �M S      E  , ,  �� Qu  �� R=  � R=  � Qu  �� Qu      E  , ,  �� S  �� S�  � S�  � S  �� S      E  , ,  �m Qu  �m R=  �5 R=  �5 Qu  �m Qu      E  , ,  �m S  �m S�  �5 S�  �5 S  �m S      E  , ,  �� Qu  �� R=  �� R=  �� Qu  �� Qu      E  , ,  �� S  �� S�  �� S�  �� S  �� S      E  , ,  � Qu  � R=  �U R=  �U Qu  � Qu      E  , ,  � S  � S�  �U S�  �U S  � S      E  , ,  � Qu  � R=  �� R=  �� Qu  � Qu      E  , ,  � S  � S�  �� S�  �� S  � S      E  , ,  � Qu  � R=  �u R=  �u Qu  � Qu      E  , ,  � S  � S�  �u S�  �u S  � S      E  , ,  �= Qu  �= R=  � R=  � Qu  �= Qu      E  , ,  �= S  �= S�  � S�  � S  �= S      E  , ,  �� Qu  �� R=  � R=  � Qu  �� Qu      E  , ,  �� S  �� S�  � S�  � S  �� S      E  , ,  �] Qu  �] R=  �% R=  �% Qu  �] Qu      E  , ,  �] S  �] S�  �% S�  �% S  �] S      E  , ,  �� Qu  �� R=  � R=  � Qu  �� Qu      E  , ,  �� S  �� S�  � S�  � S  �� S      E  , ,  �} Qu  �} R=  �E R=  �E Qu  �} Qu      E  , ,  �} S  �} S�  �E S�  �E S  �} S      E  , ,  � Qu  � R=  �� R=  �� Qu  � Qu      E  , ,  � S  � S�  �� S�  �� S  � S      E  , ,  �� Qu  �� R=  �e R=  �e Qu  �� Qu      E  , ,  �� S  �� S�  �e S�  �e S  �� S      E  , ,  �- Qu  �- R=  �� R=  �� Qu  �- Qu      E  , ,  �- S  �- S�  �� S�  �� S  �- S      E  , ,  �� Cg  �� D/  � D/  � Cg  �� Cg      E  , ,  �a Cg  �a D/  �) D/  �) Cg  �a Cg      E  , ,  �� A�  �� B�  � B�  � A�  �� A�      E  , ,  �� @G  �� A  � A  � @G  �� @G      E  , ,  �a @G  �a A  �) A  �) @G  �a @G      E  , ,  �a A�  �a B�  �) B�  �) A�  �a A�      E  , ,  �� 5W  �� 6  � 6  � 5W  �� 5W      E  , ,  �a 5W  �a 6  �) 6  �) 5W  �a 5W      E  , ,  �� 6�  �� 7�  � 7�  � 6�  �� 6�      E  , ,  �a 6�  �a 7�  �) 7�  �) 6�  �a 6�      E  , ,  �� 8w  �� 9?  � 9?  � 8w  �� 8w      E  , ,  �a 8w  �a 9?  �) 9?  �) 8w  �a 8w      E  , ,  �� :  �� :�  � :�  � :  �� :      E  , ,  �a :  �a :�  �) :�  �) :  �a :      E  , ,  �� ;�  �� <_  � <_  � ;�  �� ;�      E  , ,  �a ;�  �a <_  �) <_  �) ;�  �a ;�      E  , ,  �� ='  �� =�  � =�  � ='  �� ='      E  , ,  �a ='  �a =�  �) =�  �) ='  �a ='      E  , ,  �� >�  �� ?  � ?  � >�  �� >�      E  , ,  �a >�  �a ?  �) ?  �) >�  �a >�      E  , , N S N S� N� S� N� S N S      E  , , O� Qu O� R= Pu R= Pu Qu O� Qu      E  , , O� S O� S� Pu S� Pu S O� S      E  , , = Qu = R=   R=   Qu = Qu      E  , , = S = S�   S�   S = S      E  , ,  � Qu  � R= !� R= !� Qu  � Qu      E  , , Y S Y S� Y� S� Y� S Y S      E  , ,  � S  � S� !� S� !� S  � S      E  , , "] Qu "] R= #% R= #% Qu "] Qu      E  , , "] S "] S� #% S� #% S "] S      E  , , #� Qu #� R= $� R= $� Qu #� Qu      E  , , #� S #� S� $� S� $� S #� S      E  , , %} Qu %} R= &E R= &E Qu %} Qu      E  , , %} S %} S� &E S� &E S %} S      E  , , ' Qu ' R= '� R= '� Qu ' Qu      E  , , ' S ' S� '� S� '� S ' S      E  , , (� Qu (� R= )e R= )e Qu (� Qu      E  , , (� S (� S� )e S� )e S (� S      E  , , *- Qu *- R= *� R= *� Qu *- Qu      E  , , *- S *- S� *� S� *� S *- S      E  , , +� Qu +� R= ,� R= ,� Qu +� Qu      E  , , +� S +� S� ,� S� ,� S +� S      E  , , -M Qu -M R= . R= . Qu -M Qu      E  , , -M S -M S� . S� . S -M S      E  , , .� Qu .� R= /� R= /� Qu .� Qu      E  , , Z� Qu Z� R= [e R= [e Qu Z� Qu      E  , , Z� S Z� S� [e S� [e S Z� S      E  , , \- Qu \- R= \� R= \� Qu \- Qu      E  , , \- S \- S� \� S� \� S \- S      E  , , ]� Qu ]� R= ^� R= ^� Qu ]� Qu      E  , , ]� S ]� S� ^� S� ^� S ]� S      E  , , _M Qu _M R= ` R= ` Qu _M Qu      E  , , _M S _M S� ` S� ` S _M S      E  , , `� Qu `� R= a� R= a� Qu `� Qu      E  , , `� S `� S� a� S� a� S `� S      E  , , bm Qu bm R= c5 R= c5 Qu bm Qu      E  , , bm S bm S� c5 S� c5 S bm S      E  , , c� Qu c� R= d� R= d� Qu c� Qu      E  , , c� S c� S� d� S� d� S c� S      E  , , .� S .� S� /� S� /� S .� S      E  , , 0m Qu 0m R= 15 R= 15 Qu 0m Qu      E  , , 0m S 0m S� 15 S� 15 S 0m S      E  , , 1� Qu 1� R= 2� R= 2� Qu 1� Qu      E  , , 1� S 1� S� 2� S� 2� S 1� S      E  , , 3� Qu 3� R= 4U R= 4U Qu 3� Qu      E  , , 3� S 3� S� 4U S� 4U S 3� S      E  , , 5 Qu 5 R= 5� R= 5� Qu 5 Qu      E  , , 5 S 5 S� 5� S� 5� S 5 S      E  , , 6� Qu 6� R= 7u R= 7u Qu 6� Qu      E  , , 6� S 6� S� 7u S� 7u S 6� S      E  , , 8= Qu 8= R= 9 R= 9 Qu 8= Qu      E  , , 8= S 8= S� 9 S� 9 S 8= S      E  , , 9� Qu 9� R= :� R= :� Qu 9� Qu      E  , , 9� S 9� S� :� S� :� S 9� S      E  , , ;] Qu ;] R= <% R= <% Qu ;] Qu      E  , , Q= Qu Q= R= R R= R Qu Q= Qu      E  , , ;] S ;] S� <% S� <% S ;] S      E  , , <� Qu <� R= =� R= =� Qu <� Qu      E  , , <� S <� S� =� S� =� S <� S      E  , , >} Qu >} R= ?E R= ?E Qu >} Qu      E  , , >} S >} S� ?E S� ?E S >} S      E  , , @ Qu @ R= @� R= @� Qu @ Qu      E  , , @ S @ S� @� S� @� S @ S      E  , , A� Qu A� R= Be R= Be Qu A� Qu      E  , , A� S A� S� Be S� Be S A� S      E  , , C- Qu C- R= C� R= C� Qu C- Qu      E  , , C- S C- S� C� S� C� S C- S      E  , , D� Qu D� R= E� R= E� Qu D� Qu      E  , , D� S D� S� E� S� E� S D� S      E  , , FM Qu FM R= G R= G Qu FM Qu      E  , , FM S FM S� G S� G S FM S      E  , , G� Qu G� R= H� R= H� Qu G� Qu      E  , , G� S G� S� H� S� H� S G� S      E  , , Im Qu Im R= J5 R= J5 Qu Im Qu      E  , , Im S Im S� J5 S� J5 S Im S      E  , , J� Qu J� R= K� R= K� Qu J� Qu      E  , , Q= S Q= S� R S� R S Q= S      E  , , R� Qu R� R= S� R= S� Qu R� Qu      E  , , R� S R� S� S� S� S� S R� S      E  , , T] Qu T] R= U% R= U% Qu T] Qu      E  , , T] S T] S� U% S� U% S T] S      E  , , U� Qu U� R= V� R= V� Qu U� Qu      E  , , U� S U� S� V� S� V� S U� S      E  , , W} Qu W} R= XE R= XE Qu W} Qu      E  , , W} S W} S� XE S� XE S W} S      E  , , Y Qu Y R= Y� R= Y� Qu Y Qu      E  , , J� S J� S� K� S� K� S J� S      E  , , L� Qu L� R= MU R= MU Qu L� Qu      E  , , L� S L� S� MU S� MU S L� S      E  , , N Qu N R= N� R= N� Qu N Qu      E  , ,  �� ��  �� �o  � �o  � ��  �� ��      E  , ,  �a ��  �a �o  �) �o  �) ��  �a ��      E  , ,  ��  7  ��  �  �  �  �  7  ��  7      E  , ,  �a  7  �a  �  �)  �  �)  7  �a  7      E  , ,  �� �  �� �  � �  � �  �� �      E  , ,  �a �  �a �  �) �  �) �  �a �      E  , ,  �� W  ��   �   � W  �� W      E  , ,  �a W  �a   �)   �) W  �a W      E  , ,  �� �  �� �  � �  � �  �� �      E  , ,  �a �  �a �  �) �  �) �  �a �      E  , ,  �� w  �� ?  � ?  � w  �� w      E  , ,  �a w  �a ?  �) ?  �) w  �a w      E  , ,  ��   �� �  � �  �   ��       E  , ,  �a   �a �  �) �  �)   �a       E  , ,  �� 	�  �� 
_  � 
_  � 	�  �� 	�      E  , ,  �a 	�  �a 
_  �) 
_  �) 	�  �a 	�      E  , ,  �� '  �� �  � �  � '  �� '      E  , ,  �a '  �a �  �) �  �) '  �a '      E  , ,  �� �  ��   �   � �  �� �      E  , ,  �a �  �a   �)   �) �  �a �      E  , ,  �� G  ��   �   � G  �� G      E  , ,  �a G  �a   �)   �) G  �a G      E  , ,  �� �  �� �  � �  � �  �� �      E  , ,  �a �  �a �  �) �  �) �  �a �      E  , ,  �� g  �� /  � /  � g  �� g      E  , ,  �a g  �a /  �) /  �) g  �a g      E  , ,  �� �  �� �  � �  � �  �� �      E  , ,  �a �  �a �  �) �  �) �  �a �      E  , ,  �� �  �� O  � O  � �  �� �      E  , ,  �a �  �a O  �) O  �) �  �a �      E  , ,  ��   �� �  � �  �   ��       E  , ,  �a   �a �  �) �  �)   �a       E  , ,  �� �  �� o  � o  � �  �� �      E  , ,  �a �  �a o  �) o  �) �  �a �      E  , ,  �� 7  �� �  � �  � 7  �� 7      E  , ,  �a 7  �a �  �) �  �) 7  �a 7      E  , ,  �� �  �� �  � �  � �  �� �      E  , ,  �a �  �a �  �) �  �) �  �a �      E  , ,  �� W  ��   �   � W  �� W      E  , ,  �a W  �a   �)   �) W  �a W      E  , ,  �� �  �� �  � �  � �  �� �      E  , ,  �a �  �a �  �) �  �) �  �a �      E  , ,  �� w  ��  ?  �  ?  � w  �� w      E  , ,  �a w  �a  ?  �)  ?  �) w  �a w      E  , ,  �� !  �� !�  � !�  � !  �� !      E  , ,  �a !  �a !�  �) !�  �) !  �a !      E  , ,  �� "�  �� #_  � #_  � "�  �� "�      E  , ,  �a "�  �a #_  �) #_  �) "�  �a "�      E  , ,  �� $'  �� $�  � $�  � $'  �� $'      E  , ,  �a $'  �a $�  �) $�  �) $'  �a $'      E  , ,  �� %�  �� &  � &  � %�  �� %�      E  , ,  �a %�  �a &  �) &  �) %�  �a %�      E  , ,  �� 'G  �� (  � (  � 'G  �� 'G      E  , ,  �a 'G  �a (  �) (  �) 'G  �a 'G      E  , ,  �� (�  �� )�  � )�  � (�  �� (�      E  , ,  �a (�  �a )�  �) )�  �) (�  �a (�      E  , ,  �� *g  �� +/  � +/  � *g  �� *g      E  , ,  �a *g  �a +/  �) +/  �) *g  �a *g      E  , ,  �� +�  �� ,�  � ,�  � +�  �� +�      E  , ,  �a +�  �a ,�  �) ,�  �) +�  �a +�      E  , ,  �� -�  �� .O  � .O  � -�  �� -�      E  , ,  �a -�  �a .O  �) .O  �) -�  �a -�      E  , ,  �� /  �� /�  � /�  � /  �� /      E  , ,  �a /  �a /�  �) /�  �) /  �a /      E  , ,  �� 0�  �� 1o  � 1o  � 0�  �� 0�      E  , ,  �a 0�  �a 1o  �) 1o  �) 0�  �a 0�      E  , ,  �� 27  �� 2�  � 2�  � 27  �� 27      E  , ,  �a 27  �a 2�  �) 2�  �) 27  �a 27      E  , ,  �� �  �� �_  � �_  � �  �� �      E  , ,  �a �  �a �_  �) �_  �) �  �a �      E  , ,  �� �'  �� ��  � ��  � �'  �� �'      E  , ,  �a �'  �a ��  �) ��  �) �'  �a �'      E  , ,  �� �  �� �  � �  � �  �� �      E  , ,  �a �  �a �  �) �  �) �  �a �      E  , ,  �� �G  �� �  � �  � �G  �� �G      E  , ,  �a �G  �a �  �) �  �) �G  �a �G      E  , ,  �� �W  �� �  � �  � �W  �� �W      E  , ,  �a �W  �a �  �) �  �) �W  �a �W      E  , ,  �� ��  �� �  � �  � ��  �� ��      E  , ,  �a ��  �a �  �) �  �) ��  �a ��      E  , ,  �� ��  �� ��  � ��  � ��  �� ��      E  , ,  �a ��  �a ��  �) ��  �) ��  �a ��      E  , ,  �� �g  �� �/  � �/  � �g  �� �g      E  , ,  �a �g  �a �/  �) �/  �) �g  �a �g      E  , ,  �� ��  �� ��  � ��  � ��  �� ��      E  , ,  �a ��  �a ��  �) ��  �) ��  �a ��      E  , ,  �� ��  �� �O  � �O  � ��  �� ��      E  , ,  �a ��  �a �O  �) �O  �) ��  �a ��      E  , ,  �� �  �� ��  � ��  � �  �� �      E  , ,  �a ��  �a �  �) �  �) ��  �a ��      E  , ,  �� ��  �� ȿ  � ȿ  � ��  �� ��      E  , ,  �a ��  �a ȿ  �) ȿ  �) ��  �a ��      E  , ,  �� ɇ  �� �O  � �O  � ɇ  �� ɇ      E  , ,  �a ɇ  �a �O  �) �O  �) ɇ  �a ɇ      E  , ,  �� �  �� ��  � ��  � �  �� �      E  , ,  �a �  �a ��  �) ��  �) �  �a �      E  , ,  �� ̧  �� �o  � �o  � ̧  �� ̧      E  , ,  �a ̧  �a �o  �) �o  �) ̧  �a ̧      E  , ,  �� �7  �� ��  � ��  � �7  �� �7      E  , ,  �a �7  �a ��  �) ��  �) �7  �a �7      E  , ,  �� ��  �� Џ  � Џ  � ��  �� ��      E  , ,  �a ��  �a Џ  �) Џ  �) ��  �a ��      E  , ,  �� �W  �� �  � �  � �W  �� �W      E  , ,  �a �W  �a �  �) �  �) �W  �a �W      E  , ,  �� ��  �� ӯ  � ӯ  � ��  �� ��      E  , ,  �a ��  �a ӯ  �) ӯ  �) ��  �a ��      E  , ,  �� �w  �� �?  � �?  � �w  �� �w      E  , ,  �a �  �a ��  �) ��  �) �  �a �      E  , ,  �a ��  �a �  �) �  �) ��  �a ��      E  , ,  �� �  �� �O  � �O  � �  �� �      E  , ,  �a �  �a �O  �) �O  �) �  �a �      E  , ,  �� �  �� ��  � ��  � �  �� �      E  , ,  �a �  �a ��  �) ��  �) �  �a �      E  , ,  �� �  �� �o  � �o  � �  �� �      E  , ,  �a �  �a �o  �) �o  �) �  �a �      E  , ,  �� �7  �� ��  � ��  � �7  �� �7      E  , ,  �a �7  �a ��  �) ��  �) �7  �a �7      E  , ,  �� ��  �� �  � �  � ��  �� ��      E  , ,  �� �w  �� �?  � �?  � �w  �� �w      E  , ,  �a �w  �a �?  �) �?  �) �w  �a �w      E  , ,  �� �  �� ��  � ��  � �  �� �      E  , ,  �a �  �a ��  �) ��  �) �  �a �      E  , ,  �a �w  �a �?  �) �?  �) �w  �a �w      E  , ,  �� �  �� ��  � ��  � �  �� �      E  , ,  �a �  �a ��  �) ��  �) �  �a �      E  , ,  �� ח  �� �_  � �_  � ח  �� ח      E  , ,  �a ח  �a �_  �) �_  �) ח  �a ח      E  , ,  �� �'  �� ��  � ��  � �'  �� �'      E  , ,  �a �'  �a ��  �) ��  �) �'  �a �'      E  , ,  �� ڷ  �� �  � �  � ڷ  �� ڷ      E  , ,  �a ڷ  �a �  �) �  �) ڷ  �a ڷ      E  , ,  �� �G  �� �  � �  � �G  �� �G      E  , ,  �a �G  �a �  �) �  �) �G  �a �G      E  , ,  �� ��  �� ޟ  � ޟ  � ��  �� ��      E  , ,  �a ��  �a ޟ  �) ޟ  �) ��  �a ��      E  , ,  �� �g  �� �/  � �/  � �g  �� �g      E  , ,  �a �g  �a �/  �) �/  �) �g  �a �g      E  , ,  �� ��  �� �  � �  � ��  �� ��      E  , , � Z� � [� [ [� [ Z� � Z�      E  , ,  Z�  [� � [� � Z�  Z�      E  , , d� 3� d� 4� e� 4� e� 3� d� 3�      E  , , d� 2) d� 2� e� 2� e� 2) d� 2)      E  , ,  �a ��  �a �O  �) �O  �) ��  �a ��      E  , ,  �� �  �� ��  � ��  � �  �� �      E  , ,  �a �  �a ��  �) ��  �) �  �a �      E  , ,  �� ��  �� �o  � �o  � ��  �� ��      E  , ,  �a ��  �a �o  �) �o  �) ��  �a ��      E  , ,  �� �7  �� ��  � ��  � �7  �� �7      E  , ,  �a �7  �a ��  �) ��  �) �7  �a �7      E  , ,  �� ��  �� ��  � ��  � ��  �� ��      E  , ,  �a ��  �a ��  �) ��  �) ��  �a ��      E  , ,  �� �W  �� �  � �  � �W  �� �W      E  , ,  �a �W  �a �  �) �  �) �W  �a �W      E  , ,  �� ��  �� ��  � ��  � ��  �� ��      E  , ,  �a ��  �a ��  �) ��  �) ��  �a ��      E  , ,  �� �w  �� �?  � �?  � �w  �� �w      E  , ,  �a �w  �a �?  �) �?  �) �w  �a �w      E  , ,  �� �  �� ��  � ��  � �  �� �      E  , ,  �a �  �a ��  �) ��  �) �  �a �      E  , ,  �� ��  �� �_  � �_  � ��  �� ��      E  , ,  �a ��  �a �_  �) �_  �) ��  �a ��      E  , ,  �� �'  �� ��  � ��  � �'  �� �'      E  , ,  �a �'  �a ��  �) ��  �) �'  �a �'      E  , ,  �� ��  �� �  � �  � ��  �� ��      E  , ,  �a ��  �a �  �) �  �) ��  �a ��      E  , ,  �� �G  �� �  � �  � �G  �� �G      E  , ,  �a �G  �a �  �) �  �) �G  �a �G      E  , ,  �� ��  �� ş  � ş  � ��  �� ��      E  , ,  �a ��  �a ş  �) ş  �) ��  �a ��      E  , ,  �� �g  �� �/  � �/  � �g  �� �g      E  , ,  �a �g  �a �/  �) �/  �) �g  �a �g      E  , ,  �� �G  �� �  � �  � �G  �� �G      E  , ,  �a �G  �a �  �) �  �) �G  �a �G      E  , ,  �� ��  �� ��  � ��  � ��  �� ��      E  , ,  �a ��  �a ��  �) ��  �) ��  �a ��      E  , ,  �� �g  �� �/  � �/  � �g  �� �g      E  , ,  �a �g  �a �/  �) �/  �) �g  �a �g      E  , ,  �� ��  �� ��  � ��  � ��  �� ��      E  , , � �� � �s [ �s [ �� � ��      E  , ,  ��  �s � �s � ��  ��      E  , , � �; � � [ � [ �; � �;      E  , ,  �;  � � � � �;  �;      E  , , � �� � �� [ �� [ �� � ��      E  , ,  ��  �� � �� � ��  ��      E  , , � �[ � �# [ �# [ �[ � �[      E  , ,  �[  �# � �# � �[  �[      E  , , � �� � �� [ �� [ �� � ��      E  , ,  ��  �� � �� � ��  ��      E  , , � �{ � �C [ �C [ �{ � �{      E  , ,  �{  �C � �C � �{  �{      E  , , � � � �� [ �� [ � � �      E  , ,  �  �� � �� � �  �      E  , , � �� � �c [ �c [ �� � ��      E  , ,  ��  �c � �c � ��  ��      E  , ,  �a ��  �a ��  �) ��  �) ��  �a ��      E  , ,  �� ��  �� �O  � �O  � ��  �� ��      E  , , � �+ � �� [ �� [ �+ � �+      E  , ,  �+  �� � �� � �+  �+      E  , , � �� � �� [ �� [ �� � ��      E  , ,  ��  �� � �� � ��  ��      E  , , � �K � � [ � [ �K � �K      E  , ,  �K  � � � � �K  �K      E  , , � �� � �� [ �� [ �� � ��      E  , ,  ��  �� � �� � ��  ��      E  , , � p� � q� [ q� [ p� � p�      E  , ,  p�  q� � q� � p�  p�      E  , , � rk � s3 [ s3 [ rk � rk      E  , ,  rk  s3 � s3 � rk  rk      E  , , � s� � t� [ t� [ s� � s�      E  , ,  s�  t� � t� � s�  s�      E  , , � u� � vS [ vS [ u� � u�      E  , ,  u�  vS � vS � u�  u�      E  , , � w � w� [ w� [ w � w      E  , ,  w  w� � w� � w  w      E  , , � x� � ys [ ys [ x� � x�      E  , ,  x�  ys � ys � x�  x�      E  , , � z; � { [ { [ z; � z;      E  , ,  z;  { � { � z;  z;      E  , , � {� � |� [ |� [ {� � {�      E  , ,  {�  |� � |� � {�  {�      E  , , � }[ � ~# [ ~# [ }[ � }[      E  , ,  }[  ~# � ~# � }[  }[      E  , , � ~� � � [ � [ ~� � ~�      E  , ,  ~�  � � � � ~�  ~�      E  , , � �{ � �C [ �C [ �{ � �{      E  , ,  �{  �C � �C � �{  �{      E  , , � � � �� [ �� [ � � �      E  , ,  �  �� � �� � �  �      E  , , � �� � �c [ �c [ �� � ��      E  , ,  ��  �c � �c � ��  ��      E  , , � �+ � �� [ �� [ �+ � �+      E  , ,  �+  �� � �� � �+  �+      E  , , � �� � �� [ �� [ �� � ��      E  , ,  ��  �� � �� � ��  ��      E  , , � �K � � [ � [ �K � �K      E  , ,  �K  � � � � �K  �K      E  , , � �� � �� [ �� [ �� � ��      E  , ,  ��  �� � �� � ��  ��      E  , , � �k � �3 [ �3 [ �k � �k      E  , ,  �k  �3 � �3 � �k  �k      E  , , � �� � �� [ �� [ �� � ��      E  , ,  ��  �� � �� � ��  ��      E  , , � �� � �S [ �S [ �� � ��      E  , ,  ��  �S � �S � ��  ��      E  , , � � � �� [ �� [ � � �      E  , ,  �  �� � �� � �  �      E  , , � \� � ]S [ ]S [ \� � \�      E  , ,  \�  ]S � ]S � \�  \�      E  , , � ^ � ^� [ ^� [ ^ � ^      E  , ,  ^  ^� � ^� � ^  ^      E  , , � _� � `s [ `s [ _� � _�      E  , ,  _�  `s � `s � _�  _�      E  , , � a; � b [ b [ a; � a;      E  , ,  a;  b � b � a;  a;      E  , , � b� � c� [ c� [ b� � b�      E  , ,  b�  c� � c� � b�  b�      E  , , � d[ � e# [ e# [ d[ � d[      E  , ,  d[  e# � e# � d[  d[      E  , , � e� � f� [ f� [ e� � e�      E  , ,  e�  f� � f� � e�  e�      E  , , � g{ � hC [ hC [ g{ � g{      E  , ,  g{  hC � hC � g{  g{      E  , , � i � i� [ i� [ i � i      E  , ,  i  i� � i� � i  i      E  , , � j� � kc [ kc [ j� � j�      E  , ,  j�  kc � kc � j�  j�      E  , , � l+ � l� [ l� [ l+ � l+      E  , ,  l+  l� � l� � l+  l+      E  , , � m� � n� [ n� [ m� � m�      E  , ,  m�  n� � n� � m�  m�      E  , , � oK � p [ p [ oK � oK      E  , ,  oK  p � p � oK  oK      E  , , XY 3� XY 4� Y! 4� Y! 3� XY 3�      E  , , XY 2) XY 2� Y! 2� Y! 2) XY 2)      E  , , a� 3� a� 4� b� 4� b� 3� a� 3�      E  , , a� 2) a� 2� b� 2� b� 2) a� 2)      E  , , `) 3� `) 4� `� 4� `� 3� `) 3�      E  , , `) 2) `) 2� `� 2� `� 2) `) 2)      E  , , ^� 3� ^� 4� _a 4� _a 3� ^� 3�      E  , , ^� 2) ^� 2� _a 2� _a 2) ^� 2)      E  , , ]	 3� ]	 4� ]� 4� ]� 3� ]	 3�      E  , , ]	 2) ]	 2� ]� 2� ]� 2) ]	 2)      E  , , [y 3� [y 4� \A 4� \A 3� [y 3�      E  , , [y 2) [y 2� \A 2� \A 2) [y 2)      E  , , Y� 3� Y� 4� Z� 4� Z� 3� Y� 3�      E  , , Y� 2) Y� 2� Z� 2� Z� 2) Y� 2)      E  , , cI 3� cI 4� d 4� d 3� cI 3�      E  , , cI 2) cI 2� d 2� d 2) cI 2)      E  , , )y 3� )y 4� *A 4� *A 3� )y 3�      E  , , )y 2) )y 2� *A 2� *A 2) )y 2)      E  , , '� 3� '� 4� (� 4� (� 3� '� 3�      E  , , '� 2) '� 2� (� 2� (� 2) '� 2)      E  , , &Y 3� &Y 4� '! 4� '! 3� &Y 3�      E  , , &Y 2) &Y 2� '! 2� '! 2) &Y 2)      E  , , $� 3� $� 4� %� 4� %� 3� $� 3�      E  , , $� 2) $� 2� %� 2� %� 2) $� 2)      E  , , #9 3� #9 4� $ 4� $ 3� #9 3�      E  , , #9 2) #9 2� $ 2� $ 2) #9 2)      E  , , !� 3� !� 4� "q 4� "q 3� !� 3�      E  , , V� 3� V� 4� W� 4� W� 3� V� 3�      E  , , V� 2) V� 2� W� 2� W� 2) V� 2)      E  , , U9 3� U9 4� V 4� V 3� U9 3�      E  , , U9 2) U9 2� V 2� V 2) U9 2)      E  , , S� 3� S� 4� Tq 4� Tq 3� S� 3�      E  , , S� 2) S� 2� Tq 2� Tq 2) S� 2)      E  , , R 3� R 4� R� 4� R� 3� R 3�      E  , , R 2) R 2� R� 2� R� 2) R 2)      E  , , P� 3� P� 4� QQ 4� QQ 3� P� 3�      E  , , P� 2) P� 2� QQ 2� QQ 2) P� 2)      E  , , N� 3� N� 4� O� 4� O� 3� N� 3�      E  , , N� 2) N� 2� O� 2� O� 2) N� 2)      E  , , Mi 3� Mi 4� N1 4� N1 3� Mi 3�      E  , , Mi 2) Mi 2� N1 2� N1 2) Mi 2)      E  , , K� 3� K� 4� L� 4� L� 3� K� 3�      E  , , K� 2) K� 2� L� 2� L� 2) K� 2)      E  , , JI 3� JI 4� K 4� K 3� JI 3�      E  , , JI 2) JI 2� K 2� K 2) JI 2)      E  , , H� 3� H� 4� I� 4� I� 3� H� 3�      E  , , H� 2) H� 2� I� 2� I� 2) H� 2)      E  , , G) 3� G) 4� G� 4� G� 3� G) 3�      E  , , G) 2) G) 2� G� 2� G� 2) G) 2)      E  , , E� 3� E� 4� Fa 4� Fa 3� E� 3�      E  , , E� 2) E� 2� Fa 2� Fa 2) E� 2)      E  , , D	 3� D	 4� D� 4� D� 3� D	 3�      E  , , D	 2) D	 2� D� 2� D� 2) D	 2)      E  , , By 3� By 4� CA 4� CA 3� By 3�      E  , , By 2) By 2� CA 2� CA 2) By 2)      E  , , @� 3� @� 4� A� 4� A� 3� @� 3�      E  , , @� 2) @� 2� A� 2� A� 2) @� 2)      E  , , ?Y 3� ?Y 4� @! 4� @! 3� ?Y 3�      E  , , ?Y 2) ?Y 2� @! 2� @! 2) ?Y 2)      E  , , =� 3� =� 4� >� 4� >� 3� =� 3�      E  , , =� 2) =� 2� >� 2� >� 2) =� 2)      E  , , <9 3� <9 4� = 4� = 3� <9 3�      E  , , <9 2) <9 2� = 2� = 2) <9 2)      E  , , :� 3� :� 4� ;q 4� ;q 3� :� 3�      E  , , :� 2) :� 2� ;q 2� ;q 2) :� 2)      E  , , 9 3� 9 4� 9� 4� 9� 3� 9 3�      E  , , 9 2) 9 2� 9� 2� 9� 2) 9 2)      E  , , 7� 3� 7� 4� 8Q 4� 8Q 3� 7� 3�      E  , , 7� 2) 7� 2� 8Q 2� 8Q 2) 7� 2)      E  , , 5� 3� 5� 4� 6� 4� 6� 3� 5� 3�      E  , , 5� 2) 5� 2� 6� 2� 6� 2) 5� 2)      E  , , 4i 3� 4i 4� 51 4� 51 3� 4i 3�      E  , , 4i 2) 4i 2� 51 2� 51 2) 4i 2)      E  , , 2� 3� 2� 4� 3� 4� 3� 3� 2� 3�      E  , , 2� 2) 2� 2� 3� 2� 3� 2) 2� 2)      E  , , 1I 3� 1I 4� 2 4� 2 3� 1I 3�      E  , , 1I 2) 1I 2� 2 2� 2 2) 1I 2)      E  , , /� 3� /� 4� 0� 4� 0� 3� /� 3�      E  , , /� 2) /� 2� 0� 2� 0� 2) /� 2)      E  , , .) 3� .) 4� .� 4� .� 3� .) 3�      E  , , .) 2) .) 2� .� 2� .� 2) .) 2)      E  , , ,� 3� ,� 4� -a 4� -a 3� ,� 3�      E  , , ,� 2) ,� 2� -a 2� -a 2) ,� 2)      E  , , +	 3� +	 4� +� 4� +� 3� +	 3�      E  , , +	 2) +	 2� +� 2� +� 2) +	 2)      E  , , !� 2) !� 2� "q 2� "q 2) !� 2)      E  , ,   3�   4�  � 4�  � 3�   3�      E  , ,   2)   2�  � 2�  � 2)   2)      E  , , � 3� � 4� Q 4� Q 3� � 3�      E  , , � 2) � 2� Q 2� Q 2) � 2)      E  , , � 'k � (3 [ (3 [ 'k � 'k      E  , ,  'k  (3 � (3 � 'k  'k      E  , , � (� � )� [ )� [ (� � (�      E  , ,  (�  )� � )� � (�  (�      E  , , � *� � +S [ +S [ *� � *�      E  , ,  *�  +S � +S � *�  *�      E  , ,  L�  M� � M� � L�  L�      E  , , � N{ � OC [ OC [ N{ � N{      E  , , � , � ,� [ ,� [ , � ,      E  , ,  ,  ,� � ,� � ,  ,      E  , , � -� � .s [ .s [ -� � -�      E  , ,  -�  .s � .s � -�  -�      E  , , � /; � 0 [ 0 [ /; � /;      E  , ,  /;  0 � 0 � /;  /;      E  , , � 0� � 1� [ 1� [ 0� � 0�      E  , ,  0�  1� � 1� � 0�  0�      E  , , � 2[ � 3# [ 3# [ 2[ � 2[      E  , ,  2[  3# � 3# � 2[  2[      E  , , � 3� � 4� [ 4� [ 3� � 3�      E  , ,  3�  4� � 4� � 3�  3�      E  , , � 5{ � 6C [ 6C [ 5{ � 5{      E  , ,  5{  6C � 6C � 5{  5{      E  , , � 7 � 7� [ 7� [ 7 � 7      E  , ,  7  7� � 7� � 7  7      E  , , � 8� � 9c [ 9c [ 8� � 8�      E  , ,  8�  9c � 9c � 8�  8�      E  , , � VK � W [ W [ VK � VK      E  , ,  VK  W � W � VK  VK      E  , , � W� � X� [ X� [ W� � W�      E  , ,  W�  X� � X� � W�  W�      E  , , � Yk � Z3 [ Z3 [ Yk � Yk      E  , ,  Yk  Z3 � Z3 � Yk  Yk      E  , , � :+ � :� [ :� [ :+ � :+      E  , , � L� � M� [ M� [ L� � L�      E  , , ) 3� ) 4� � 4� � 3� ) 3�      E  , , ) 2) ) 2� � 2� � 2) ) 2)      E  , , � 3� � 4� a 4� a 3� � 3�      E  , , � 2) � 2� a 2� a 2) � 2)      E  , , 	 3� 	 4� � 4� � 3� 	 3�      E  , , 	 2) 	 2� � 2� � 2) 	 2)      E  , , y 3� y 4� A 4� A 3� y 3�      E  , , y 2) y 2� A 2� A 2) y 2)      E  , , � 3� � 4� � 4� � 3� � 3�      E  , , � 2) � 2� � 2� � 2) � 2)      E  , , Y 3� Y 4� ! 4� ! 3� Y 3�      E  , , Y 2) Y 2� ! 2� ! 2) Y 2)      E  , , � 3� � 4� � 4� � 3� � 3�      E  , , � 2) � 2� � 2� � 2) � 2)      E  , ,  T�  U� � U� � T�  T�      E  , , � I� � J� [ J� [ I� � I�      E  , ,  I�  J� � J� � I�  I�      E  , , � K[ � L# [ L# [ K[ � K[      E  , ,  K[  L# � L# � K[  K[      E  , ,  H;  I � I � H;  H;      E  , , � %� � &� [ &� [ %� � %�      E  , ,  %�  &� � &� � %�  %�      E  , , � 3� � 4� � 4� � 3� � 3�      E  , , � 2) � 2� � 2� � 2) � 2)      E  , , i 3� i 4� 1 4� 1 3� i 3�      E  , , i 2) i 2� 1 2� 1 2) i 2)      E  , , � 3� � 4� � 4� � 3� � 3�      E  , , � 2) � 2� � 2� � 2) � 2)      E  , , I 3� I 4�  4�  3� I 3�      E  , , I 2) I 2�  2�  2) I 2)      E  , , � 3� � 4� � 4� � 3� � 3�      E  , , � 2) � 2� � 2� � 2) � 2)      E  , ,  N{  OC � OC � N{  N{      E  , , � P � P� [ P� [ P � P      E  , ,  P  P� � P� � P  P      E  , , � Q� � Rc [ Rc [ Q� � Q�      E  , ,  Q�  Rc � Rc � Q�  Q�      E  , , � S+ � S� [ S� [ S+ � S+      E  , ,  S+  S� � S� � S+  S+      E  , , � T� � U� [ U� [ T� � T�      E  , ,  :+  :� � :� � :+  :+      E  , , � ;� � <� [ <� [ ;� � ;�      E  , ,  ;�  <� � <� � ;�  ;�      E  , , � =K � > [ > [ =K � =K      E  , ,  =K  > � > � =K  =K      E  , , � >� � ?� [ ?� [ >� � >�      E  , ,  >�  ?� � ?� � >�  >�      E  , , � @k � A3 [ A3 [ @k � @k      E  , ,  @k  A3 � A3 � @k  @k      E  , , � A� � B� [ B� [ A� � A�      E  , ,  A�  B� � B� � A�  A�      E  , , � C� � DS [ DS [ C� � C�      E  , ,  C�  DS � DS � C�  C�      E  , , � E � E� [ E� [ E � E      E  , ,  E  E� � E� � E  E      E  , , � F� � Gs [ Gs [ F� � F�      E  , ,  F�  Gs � Gs � F�  F�      E  , , � H; � I [ I [ H; � H;      E  , , � k � 3 [ 3 [ k � k      E  , ,  k  3 � 3 � k  k      E  , , � � � � [ � [ � � �      E  , ,  �  � � � � �  �      E  , , � � � S [ S [ � � �      E  , ,  �  S � S � �  �      E  , , �  � � [ � [  �       E  , ,    � � � �         E  , , � � � s [ s [ � � �      E  , ,  �  s � s � �  �      E  , , � ; �  [  [ ; � ;      E  , ,  ;   �  � ;  ;      E  , , � � � � [ � [ � � �      E  , ,  �  � � � � �  �      E  , , � [ � # [ # [ [ � [      E  , ,  [  # � # � [  [      E  , , � { � C [ C [ { � {      E  , ,  {  C � C � {  {      E  , , �  � � [ � [  �       E  , ,    � � � �         E  , , � � �  c [  c [ � � �      E  , ,  �   c �  c � �  �      E  , , � !+ � !� [ !� [ !+ � !+      E  , ,  !+  !� � !� � !+  !+      E  , , � "� � #� [ #� [ "� � "�      E  , ,  "�  #� � #� � "�  "�      E  , , � $K � % [ % [ $K � $K      E  , ,  $K  % � % � $K  $K      E  , , � 	� � 
� [ 
� [ 	� � 	�      E  , ,  	�  
� � 
� � 	�  	�      E  , , � K �  [  [ K � K      E  , ,  K   �  � K  K      E  , , � � � � [ � [ � � �      E  , ,  �  � � � � �  �      E  , , � � � � [ � [ � � �      E  , ,  �  � � � � �  �      E  , , �� Y2 �� Y� �� Y� �� Y2 �� Y2      E  , , �� W� �� Xj �� Xj �� W� �� W�      E  , , �� W� �� Xj �� Xj �� W� �� W�      E  , , �l Y2 �l Y� �4 Y� �4 Y2 �l Y2      E  , , �l W� �l Xj �4 Xj �4 W� �l W�      E  , , �� Y2 �� Y� �� Y� �� Y2 �� Y2      E  , , �� W� �� Xj �� Xj �� W� �� W�      E  , , �L Y2 �L Y� � Y� � Y2 �L Y2      E  , , �L W� �L Xj � Xj � W� �L W�      E  , , �� Y2 �� Y� �� Y� �� Y2 �� Y2      E  , , �� W� �� Xj �� Xj �� W� �� W�      E  , , �, Y2 �, Y� �� Y� �� Y2 �, Y2      E  , , �, W� �, Xj �� Xj �� W� �, W�      E  , , �� Y2 �� Y� �d Y� �d Y2 �� Y2      E  , , �� W� �� Xj �d Xj �d W� �� W�      E  , , � Y2 � Y� �� Y� �� Y2 � Y2      E  , , � W� � Xj �� Xj �� W� � W�      E  , , �| Y2 �| Y� �D Y� �D Y2 �| Y2      E  , , �| W� �| Xj �D Xj �D W� �| W�      E  , , �� W� �� Xj �T Xj �T W� �� W�      E  , , �� Y2 �� Y� �� Y� �� Y2 �� Y2      E  , , ɜ W� ɜ Xj �d Xj �d W� ɜ W�      E  , , � Y2 � Y� �� Y� �� Y2 � Y2      E  , , � W� � Xj �� Xj �� W� � W�      E  , , �| Y2 �| Y� �D Y� �D Y2 �| Y2      E  , , �| W� �| Xj �D Xj �D W� �| W�      E  , , �� Y2 �� Y� Ŵ Y� Ŵ Y2 �� Y2      E  , , �� W� �� Xj Ŵ Xj Ŵ W� �� W�      E  , , �\ Y2 �\ Y� �$ Y� �$ Y2 �\ Y2      E  , , �\ W� �\ Xj �$ Xj �$ W� �\ W�      E  , , �� Y2 �� Y�  Y�  Y2 �� Y2      E  , , �� W� �� Xj  Xj  W� �� W�      E  , , �< Y2 �< Y� � Y� � Y2 �< Y2      E  , , �< W� �< Xj � Xj � W� �< W�      E  , , �� Y2 �� Y� �t Y� �t Y2 �� Y2      E  , , �� W� �� Xj �t Xj �t W� �� W�      E  , , � Y2 � Y� �� Y� �� Y2 � Y2      E  , , � Y2 � Y� �t Y� �t Y2 � Y2      E  , , � W� � Xj �t Xj �t W� � W�      E  , , � Y2 � Y� �� Y� �� Y2 � Y2      E  , , � W� � Xj �� Xj �� W� � W�      E  , , � Y2 � Y� �T Y� �T Y2 � Y2      E  , , � W� � Xj �T Xj �T W� � W�      E  , , �� Y2 �� Y� �� Y� �� Y2 �� Y2      E  , , �� W� �� Xj �� Xj �� W� �� W�      E  , , �l Y2 �l Y� �4 Y� �4 Y2 �l Y2      E  , , �l W� �l Xj �4 Xj �4 W� �l W�      E  , , �� Y2 �� Y� � Y� � Y2 �� Y2      E  , , �� W� �� Xj � Xj � W� �� W�      E  , , �L Y2 �L Y� � Y� � Y2 �L Y2      E  , , �L W� �L Xj � Xj � W� �L W�      E  , , � Y2 � Y� � Y� � Y2 � Y2      E  , , � W� � Xj � Xj � W� � W�      E  , , �, Y2 �, Y� �� Y� �� Y2 �, Y2      E  , , �, W� �, Xj �� Xj �� W� �, W�      E  , , � Y2 � Y� �d Y� �d Y2 � Y2      E  , , � W� � Xj �d Xj �d W� � W�      E  , , � Y2 � Y� �� Y� �� Y2 � Y2      E  , , � W� � Xj �� Xj �� W� � W�      E  , , �| Y2 �| Y� �D Y� �D Y2 �| Y2      E  , , �| W� �| Xj �D Xj �D W� �| W�      E  , , �� Y2 �� Y� ޴ Y� ޴ Y2 �� Y2      E  , , �� W� �� Xj ޴ Xj ޴ W� �� W�      E  , , �\ Y2 �\ Y� �$ Y� �$ Y2 �\ Y2      E  , , �\ W� �\ Xj �$ Xj �$ W� �\ W�      E  , , �� Y2 �� Y� ۔ Y� ۔ Y2 �� Y2      E  , , �� W� �� Xj ۔ Xj ۔ W� �� W�      E  , , �< Y2 �< Y� � Y� � Y2 �< Y2      E  , , �< W� �< Xj � Xj � W� �< W�      E  , , ׬ Y2 ׬ Y� �t Y� �t Y2 ׬ Y2      E  , , ׬ W� ׬ Xj �t Xj �t W� ׬ W�      E  , , � Y2 � Y� �� Y� �� Y2 � Y2      E  , , � W� � Xj �� Xj �� W� � W�      E  , , Ԍ Y2 Ԍ Y� �T Y� �T Y2 Ԍ Y2      E  , , Ԍ W� Ԍ Xj �T Xj �T W� Ԍ W�      E  , , �� Y2 �� Y� �� Y� �� Y2 �� Y2      E  , , �� W� �� Xj �� Xj �� W� �� W�      E  , , �l Y2 �l Y� �4 Y� �4 Y2 �l Y2      E  , , �l W� �l Xj �4 Xj �4 W� �l W�      E  , , �� Y2 �� Y� Ф Y� Ф Y2 �� Y2      E  , , �� W� �� Xj Ф Xj Ф W� �� W�      E  , , �L Y2 �L Y� � Y� � Y2 �L Y2      E  , , �L W� �L Xj � Xj � W� �L W�      E  , , ̼ Y2 ̼ Y� ̈́ Y� ̈́ Y2 ̼ Y2      E  , , ̼ W� ̼ Xj ̈́ Xj ̈́ W� ̼ W�      E  , , �, Y2 �, Y� �� Y� �� Y2 �, Y2      E  , , �, W� �, Xj �� Xj �� W� �, W�      E  , , ɜ Y2 ɜ Y� �d Y� �d Y2 ɜ Y2      E  , , � W� � Xj �� Xj �� W� � W�      E  , , �� Y2 �� Y� �T Y� �T Y2 �� Y2      E  , , v	 2) v	 2� v� 2� v� 2) v	 2)      E  , , ty 3� ty 4� uA 4� uA 3� ty 3�      E  , , |I 2) |I 2� } 2� } 2) |I 2)      E  , , �\ Y2 �\ Y� �$ Y� �$ Y2 �\ Y2      E  , , �\ W� �\ Xj �$ Xj �$ W� �\ W�      E  , , �� Y2 �� Y� �� Y� �� Y2 �� Y2      E  , , �� W� �� Xj �� Xj �� W� �� W�      E  , , z� 3� z� 4� {� 4� {� 3� z� 3�      E  , , z� 2) z� 2� {� 2� {� 2) z� 2)      E  , , y) 3� y) 4� y� 4� y� 3� y) 3�      E  , , y) 2) y) 2� y� 2� y� 2) y) 2)      E  , , w� 3� w� 4� xa 4� xa 3� w� 3�      E  , , fi 2) fi 2� g1 2� g1 2) fi 2)      E  , , �� 3� �� 4� �� 4� �� 3� �� 3�      E  , , �� 2) �� 2� �� 2� �� 2) �� 2)      E  , , �Y 3� �Y 4� �! 4� �! 3� �Y 3�      E  , , �Y 2) �Y 2� �! 2� �! 2) �Y 2)      E  , , �� 3� �� 4� �� 4� �� 3� �� 3�      E  , , �� 2) �� 2� �� 2� �� 2) �� 2)      E  , , �9 3� �9 4� � 4� � 3� �9 3�      E  , , �9 2) �9 2� � 2� � 2) �9 2)      E  , , �� 3� �� 4� �q 4� �q 3� �� 3�      E  , , �� 2) �� 2� �q 2� �q 2) �� 2)      E  , , � 3� � 4� �� 4� �� 3� � 3�      E  , , � 2) � 2� �� 2� �� 2) � 2)      E  , , �� 3� �� 4� �Q 4� �Q 3� �� 3�      E  , , �� 2) �� 2� �Q 2� �Q 2) �� 2)      E  , , �� 3� �� 4� �� 4� �� 3� �� 3�      E  , , �� 2) �� 2� �� 2� �� 2) �� 2)      E  , , �i 3� �i 4� �1 4� �1 3� �i 3�      E  , , �i 2) �i 2� �1 2� �1 2) �i 2)      E  , , �� 3� �� 4� �� 4� �� 3� �� 3�      E  , , �� 2) �� 2� �� 2� �� 2) �� 2)      E  , , �I 3� �I 4� � 4� � 3� �I 3�      E  , , �I 2) �I 2� � 2� � 2) �I 2)      E  , , ty 2) ty 2� uA 2� uA 2) ty 2)      E  , , w� 2) w� 2� xa 2� xa 2) w� 2)      E  , , v	 3� v	 4� v� 4� v� 3� v	 3�      E  , , r� 3� r� 4� s� 4� s� 3� r� 3�      E  , , r� 2) r� 2� s� 2� s� 2) r� 2)      E  , , qY 3� qY 4� r! 4� r! 3� qY 3�      E  , , qY 2) qY 2� r! 2� r! 2) qY 2)      E  , , o� 3� o� 4� p� 4� p� 3� o� 3�      E  , , o� 2) o� 2� p� 2� p� 2) o� 2)      E  , , n9 3� n9 4� o 4� o 3� n9 3�      E  , , n9 2) n9 2� o 2� o 2) n9 2)      E  , , l� 3� l� 4� mq 4� mq 3� l� 3�      E  , , l� 2) l� 2� mq 2� mq 2) l� 2)      E  , , k 3� k 4� k� 4� k� 3� k 3�      E  , , k 2) k 2� k� 2� k� 2) k 2)      E  , , i� 3� i� 4� jQ 4� jQ 3� i� 3�      E  , , i� 2) i� 2� jQ 2� jQ 2) i� 2)      E  , , g� 3� g� 4� h� 4� h� 3� g� 3�      E  , , g� 2) g� 2� h� 2� h� 2) g� 2)      E  , , fi 3� fi 4� g1 4� g1 3� fi 3�      E  , , �� 3� �� 4� �� 4� �� 3� �� 3�      E  , , �� 2) �� 2� �� 2� �� 2) �� 2)      E  , , �) 3� �) 4� �� 4� �� 3� �) 3�      E  , , �) 2) �) 2� �� 2� �� 2) �) 2)      E  , , �� 3� �� 4� �a 4� �a 3� �� 3�      E  , , �� 2) �� 2� �a 2� �a 2) �� 2)      E  , , �	 3� �	 4� �� 4� �� 3� �	 3�      E  , , �	 2) �	 2� �� 2� �� 2) �	 2)      E  , , �y 3� �y 4� �A 4� �A 3� �y 3�      E  , , �y 2) �y 2� �A 2� �A 2) �y 2)      E  , , �� 3� �� 4� �� 4� �� 3� �� 3�      E  , , �� 2) �� 2� �� 2� �� 2) �� 2)      E  , , �Y 3� �Y 4� �! 4� �! 3� �Y 3�      E  , , �Y 2) �Y 2� �! 2� �! 2) �Y 2)      E  , , �� 3� �� 4� �� 4� �� 3� �� 3�      E  , , �� 2) �� 2� �� 2� �� 2) �� 2)      E  , , �9 3� �9 4� � 4� � 3� �9 3�      E  , , �9 2) �9 2� � 2� � 2) �9 2)      E  , , �� 3� �� 4� �q 4� �q 3� �� 3�      E  , , �� 2) �� 2� �q 2� �q 2) �� 2)      E  , , � 3� � 4� �� 4� �� 3� � 3�      E  , , � 2) � 2� �� 2� �� 2) � 2)      E  , , �� 3� �� 4� �Q 4� �Q 3� �� 3�      E  , , �� 2) �� 2� �Q 2� �Q 2) �� 2)      E  , , �� 3� �� 4� �� 4� �� 3� �� 3�      E  , , �� 2) �� 2� �� 2� �� 2) �� 2)      E  , , i 3� i 4� �1 4� �1 3� i 3�      E  , , i 2) i 2� �1 2� �1 2) i 2)      E  , , }� 3� }� 4� ~� 4� ~� 3� }� 3�      E  , , }� 2) }� 2� ~� 2� ~� 2) }� 2)      E  , , |I 3� |I 4� } 4� } 3� |I 3�      E  , , � Z� � [~ [ [~ [ Z� � Z�      E  , , 
s Z� 
s [~ ; [~ ; Z� 
s Z�      E  , , � Z� � [~ 	� [~ 	� Z� � Z�      E  , ,  Z�  [~ � [~ � Z�  Z�      E  , , 
s �f 
s �. ; �. ; �f 
s �f      E  , , � �f � �. 	� �. 	� �f � �f      E  , ,  �f  �. � �. � �f  �f      E  , , � �f � �. [ �. [ �f � �f      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , ,  ��  �� � �� � ��  ��      E  , , � �� � �� 	� �� 	� �� � ��      E  , , � �� � �� [ �� [ �� � ��      E  , ,  �6  �� � �� � �6  �6      E  , , 
s �f 
s �. ; �. ; �f 
s �f      E  , ,  �V  � � � � �V  �V      E  , ,  ��  �n � �n � ��  ��      E  , , 
s �� 
s �^ ; �^ ; �� 
s ��      E  , ,  �  �� � �� � �  �      E  , ,  ��  �N � �N � ��  ��      E  , ,  ��  �� � �� � ��  ��      E  , , 
s � 
s �� ; �� ; � 
s �      E  , , 
s �� 
s  ;  ; �� 
s ��      E  , , � Ɔ � �N 	� �N 	� Ɔ � Ɔ      E  , , 
s �v 
s �> ; �> ; �v 
s �v      E  , , � �� � ž 	� ž 	� �� � ��      E  , ,  Ɔ  �N � �N � Ɔ  Ɔ      E  , , � �f � �. 	� �. 	� �f � �f      E  , ,  ��  ž � ž � ��  ��      E  , , � Ɔ � �N [ �N [ Ɔ � Ɔ      E  , , � �� �  	�  	� �� � ��      E  , , � �� � ž [ ž [ �� � ��      E  , , � �F � � 	� � 	� �F � �F      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , ,  �f  �. � �. � �f  �f      E  , , � �f � �. [ �. [ �f � �f      E  , , � �� � �~ 	� �~ 	� �� � ��      E  , ,  ��   �  � ��  ��      E  , , � �� �  [  [ �� � ��      E  , , � �& � �� 	� �� 	� �& � �&      E  , , � �F � � [ � [ �F � �F      E  , , � �� � �^ 	� �^ 	� �� � ��      E  , , 
s �V 
s � ; � ; �V 
s �V      E  , ,  �F  � � � � �F  �F      E  , , � �� � �~ [ �~ [ �� � ��      E  , , 
s �F 
s � ; � ; �F 
s �F      E  , , � � � �� 	� �� 	� � � �      E  , ,  ��  �~ � �~ � ��  ��      E  , , � �& � �� [ �� [ �& � �&      E  , , � �v � �> 	� �> 	� �v � �v      E  , , � �� � �^ [ �^ [ �� � ��      E  , , � �� � �� 	� �� 	� �� � ��      E  , , 
s �� 
s ž ; ž ; �� 
s ��      E  , ,  �&  �� � �� � �&  �&      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , , � � � �� [ �� [ � � �      E  , , � �V � � 	� � 	� �V � �V      E  , , � �v � �> [ �> [ �v � �v      E  , ,  ��  �^ � �^ � ��  ��      E  , , � �� � �� 	� �� 	� �� � ��      E  , , � �� � �� [ �� [ �� � ��      E  , , � �6 � �� 	� �� 	� �6 � �6      E  , , � �V � � [ � [ �V � �V      E  , , � �� � �n 	� �n 	� �� � ��      E  , ,  �  �� � �� � �  �      E  , , � �� � �� [ �� [ �� � ��      E  , , � � � �� 	� �� 	� � � �      E  , , 
s �6 
s �� ; �� ; �6 
s �6      E  , , � �6 � �� [ �� [ �6 � �6      E  , , � �� � �N 	� �N 	� �� � ��      E  , , 
s �� 
s �~ ; �~ ; �� 
s ��      E  , , 
s � 
s �� ; �� ; � 
s �      E  , , � �� � �n [ �n [ �� � ��      E  , ,  �v  �> � �> � �v  �v      E  , , 
s Ɔ 
s �N ; �N ; Ɔ 
s Ɔ      E  , , � � � �� [ �� [ � � �      E  , , 
s �� 
s �n ; �n ; �� 
s ��      E  , , � �� � �N [ �N [ �� � ��      E  , ,  ��  �� � �� � ��  ��      E  , , 
s �� 
s �N ; �N ; �� 
s ��      E  , , 
s �& 
s �� ; �� ; �& 
s �&      E  , ,  ��  �~ � �~ � ��  ��      E  , , � �F � � [ � [ �F � �F      E  , , � �& � �� [ �� [ �& � �&      E  , , 
s �V 
s � ; � ; �V 
s �V      E  , ,  ��  �� � �� � ��  ��      E  , , 
s �� 
s �^ ; �^ ; �� 
s ��      E  , , � �6 � �� [ �� [ �6 � �6      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , ,  �&  �� � �� � �&  �&      E  , , � � � �� [ �� [ � � �      E  , ,  �6  �� � �� � �6  �6      E  , , � �� � �� 	� �� 	� �� � ��      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , , � �� � �� [ �� [ �� � ��      E  , , � �� � �� [ �� [ �� � ��      E  , , 
s �F 
s � ; � ; �F 
s �F      E  , , � �� � �^ 	� �^ 	� �� � ��      E  , , � �� � �N 	� �N 	� �� � ��      E  , ,  ��  �n � �n � ��  ��      E  , ,  �f  �. � �. � �f  �f      E  , ,  ��  �^ � �^ � ��  ��      E  , , � �& � �� 	� �� 	� �& � �&      E  , , 
s �6 
s �� ; �� ; �6 
s �6      E  , ,  �  �� � �� � �  �      E  , , 
s � 
s �� ; �� ; � 
s �      E  , , � �v � �> 	� �> 	� �v � �v      E  , , � �� � �� [ �� [ �� � ��      E  , , � � � �� [ �� [ � � �      E  , ,  ��  �N � �N � ��  ��      E  , , 
s �� 
s �~ ; �~ ; �� 
s ��      E  , , � �� � �N [ �N [ �� � ��      E  , ,  ��  �� � �� � ��  ��      E  , ,  ��  �� � �� � ��  ��      E  , , 
s �� 
s �n ; �n ; �� 
s ��      E  , ,  �  �� � �� � �  �      E  , , � �� � �^ [ �^ [ �� � ��      E  , , � �6 � �� 	� �� 	� �6 � �6      E  , , � � � �� 	� �� 	� � � �      E  , , � � � �� 	� �� 	� � � �      E  , , 
s �v 
s �> ; �> ; �v 
s �v      E  , ,  �v  �> � �> � �v  �v      E  , , � �V � � 	� � 	� �V � �V      E  , , � �V � � [ � [ �V � �V      E  , ,  �F  � � � � �F  �F      E  , , 
s � 
s �� ; �� ; � 
s �      E  , , � �� � �n [ �n [ �� � ��      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , , � �� � �� [ �� [ �� � ��      E  , , � �� � �� 	� �� 	� �� � ��      E  , , � �� � �� 	� �� 	� �� � ��      E  , ,  ��  �� � �� � ��  ��      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , , � �f � �. 	� �. 	� �f � �f      E  , , 
s �& 
s �� ; �� ; �& 
s �&      E  , , � �� � �n 	� �n 	� �� � ��      E  , , 
s �� 
s �N ; �N ; �� 
s ��      E  , , � �� � �� 	� �� 	� �� � ��      E  , , 
s �f 
s �. ; �. ; �f 
s �f      E  , , � �� � �~ 	� �~ 	� �� � ��      E  , , � �F � � 	� � 	� �F � �F      E  , , � �� � �~ [ �~ [ �� � ��      E  , ,  �V  � � � � �V  �V      E  , , � �v � �> [ �> [ �v � �v      E  , , � �f � �. [ �. [ �f � �f      E  , , 
s v� 
s w� ; w� ; v� 
s v�      E  , , � } � }� 	� }� 	� } � }      E  , , � �� � �� [ �� [ �� � ��      E  , ,  �  �� � �� � �  �      E  , , � xf � y. 	� y. 	� xf � xf      E  , , � �F � � [ � [ �F � �F      E  , , � �� � �~ 	� �~ 	� �� � ��      E  , , � � � �� 	� �� 	� � � �      E  , , � �V � � [ � [ �V � �V      E  , , 
s �� 
s �~ ; �~ ; �� 
s ��      E  , ,  ��  �~ � �~ � ��  ��      E  , ,  ~�  n � n � ~�  ~�      E  , , 
s �V 
s � ; � ; �V 
s �V      E  , , � �F � � 	� � 	� �F � �F      E  , , � ~� � n 	� n 	� ~� � ~�      E  , , � {� � |N [ |N [ {� � {�      E  , , 
s �� 
s �^ ; �^ ; �� 
s ��      E  , , � v� � w� 	� w� 	� v� � v�      E  , , � v� � w� [ w� [ v� � v�      E  , ,  �v  �> � �> � �v  �v      E  , , � �� � �^ [ �^ [ �� � ��      E  , ,  v�  w� � w� � v�  v�      E  , ,  �F  � � � � �F  �F      E  , ,  �&  �� � �� � �&  �&      E  , , � �� � �� [ �� [ �� � ��      E  , ,  ��  �� � �� � ��  ��      E  , ,  ��  �� � �� � ��  ��      E  , , 
s ~� 
s n ; n ; ~� 
s ~�      E  , , � �6 � �� 	� �� 	� �6 � �6      E  , , 
s �6 
s �� ; �� ; �6 
s �6      E  , , � �� � �� [ �� [ �� � ��      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , , � y� � z� [ z� [ y� � y�      E  , ,  }  }� � }� � }  }      E  , ,  y�  z� � z� � y�  y�      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , , � �� � �^ 	� �^ 	� �� � ��      E  , , � �& � �� 	� �� 	� �& � �&      E  , ,  �6  �� � �� � �6  �6      E  , , � } � }� [ }� [ } � }      E  , ,  ��  �^ � �^ � ��  ��      E  , , � �� � �� 	� �� 	� �� � ��      E  , , 
s } 
s }� ; }� ; } 
s }      E  , ,  ��  �� � �� � ��  ��      E  , , � �� � �� 	� �� 	� �� � ��      E  , , 
s � 
s �� ; �� ; � 
s �      E  , , � �6 � �� [ �� [ �6 � �6      E  , , 
s {� 
s |N ; |N ; {� 
s {�      E  , , � �& � �� [ �� [ �& � �&      E  , ,  xf  y. � y. � xf  xf      E  , , � {� � |N 	� |N 	� {� � {�      E  , , � � � �� [ �� [ � � �      E  , , 
s �& 
s �� ; �� ; �& 
s �&      E  , , � �V � � 	� � 	� �V � �V      E  , , 
s �F 
s � ; � ; �F 
s �F      E  , , 
s y� 
s z� ; z� ; y� 
s y�      E  , ,  �V  � � � � �V  �V      E  , , 
s �v 
s �> ; �> ; �v 
s �v      E  , , � ~� � n [ n [ ~� � ~�      E  , , � y� � z� 	� z� 	� y� � y�      E  , , 
s xf 
s y. ; y. ; xf 
s xf      E  , , � �v � �> 	� �> 	� �v � �v      E  , , � �� � �~ [ �~ [ �� � ��      E  , ,  {�  |N � |N � {�  {�      E  , , � �v � �> [ �> [ �v � �v      E  , , � xf � y. [ y. [ xf � xf      E  , , 
s �� 
s �� ; �� ; �� 
s ��      E  , , � �� � �� 	� �� 	� �� � ��      E  , , 
s r& 
s r� ; r� ; r& 
s r&      E  , ,  p�  q^ � q^ � p�  p�      E  , , � h� � i� 	� i� 	� h� � h�      E  , , � _f � `. [ `. [ _f � _f      E  , , � g6 � g� [ g� [ g6 � g6      E  , , � ]� � ^� 	� ^� 	� ]� � ]�      E  , , � o � o� [ o� [ o � o      E  , , 
s g6 
s g� ; g� ; g6 
s g6      E  , , � uF � v 	� v 	� uF � uF      E  , , 
s k� 
s l� ; l� ; k� 
s k�      E  , ,  uF  v � v � uF  uF      E  , ,  `�  a� � a� � `�  `�      E  , ,  r&  r� � r� � r&  r&      E  , ,  d  d� � d� � d  d      E  , , � ]� � ^� [ ^� [ ]� � ]�      E  , , 
s p� 
s q^ ; q^ ; p� 
s p�      E  , , � r& � r� [ r� [ r& � r&      E  , ,  \F  ] � ] � \F  \F      E  , , � mv � n> 	� n> 	� mv � mv      E  , ,  h�  i� � i� � h�  h�      E  , ,  mv  n> � n> � mv  mv      E  , ,  e�  fn � fn � e�  e�      E  , ,  b�  cN � cN � b�  b�      E  , , 
s ]� 
s ^� ; ^� ; ]� 
s ]�      E  , ,  ]�  ^� � ^� � ]�  ]�      E  , , � jV � k 	� k 	� jV � jV      E  , , 
s uF 
s v ; v ; uF 
s uF      E  , , � _f � `. 	� `. 	� _f � _f      E  , , � d � d� 	� d� 	� d � d      E  , , � o � o� 	� o� 	� o � o      E  , ,  s�  t~ � t~ � s�  s�      E  , ,  g6  g� � g� � g6  g6      E  , , 
s s� 
s t~ ; t~ ; s� 
s s�      E  , ,  o  o� � o� � o  o      E  , , � p� � q^ [ q^ [ p� � p�      E  , , � g6 � g� 	� g� 	� g6 � g6      E  , , 
s o 
s o� ; o� ; o 
s o      E  , , 
s h� 
s i� ; i� ; h� 
s h�      E  , , � s� � t~ [ t~ [ s� � s�      E  , , � e� � fn [ fn [ e� � e�      E  , , � uF � v [ v [ uF � uF      E  , , 
s mv 
s n> ; n> ; mv 
s mv      E  , , 
s \F 
s ] ; ] ; \F 
s \F      E  , , � b� � cN [ cN [ b� � b�      E  , , � \F � ] [ ] [ \F � \F      E  , , � p� � q^ 	� q^ 	� p� � p�      E  , , � e� � fn 	� fn 	� e� � e�      E  , , � k� � l� [ l� [ k� � k�      E  , , 
s jV 
s k ; k ; jV 
s jV      E  , , 
s _f 
s `. ; `. ; _f 
s _f      E  , ,  _f  `. � `. � _f  _f      E  , , � s� � t~ 	� t~ 	� s� � s�      E  , ,  jV  k � k � jV  jV      E  , , 
s d 
s d� ; d� ; d 
s d      E  , , 
s e� 
s fn ; fn ; e� 
s e�      E  , , � b� � cN 	� cN 	� b� � b�      E  , , � h� � i� [ i� [ h� � h�      E  , , � `� � a� [ a� [ `� � `�      E  , ,  k�  l� � l� � k�  k�      E  , , 
s `� 
s a� ; a� ; `� 
s `�      E  , , � r& � r� 	� r� 	� r& � r&      E  , , � \F � ] 	� ] 	� \F � \F      E  , , � k� � l� 	� l� 	� k� � k�      E  , , � jV � k [ k [ jV � jV      E  , , � `� � a� 	� a� 	� `� � `�      E  , , � d � d� [ d� [ d � d      E  , , 
s b� 
s cN ; cN ; b� 
s b�      E  , , � mv � n> [ n> [ mv � mv      E  , , -V �y -V �A . �A . �y -V �y      E  , , -V �) -V �� . �� . �) -V �)      E  , , .� �� .� �Q /� �Q /� �� .� ��      E  , , .� �� .� �� /� �� /� �� .� ��      E  , , -V �� -V �Q . �Q . �� -V ��      E  , , .� � .� �� /� �� /� � .� �      E  , , .� �	 .� �� /� �� /� �	 .� �	      E  , , -V � -V �� . �� . � -V �      E  , , .� �9 .� � /� � /� �9 .� �9      E  , , -V �9 -V � . � . �9 -V �9      E  , , .� �� .� đ /� đ /� �� .� ��      E  , , -V �� -V �� . �� . �� -V ��      E  , , -V �� -V đ . đ . �� -V ��      E  , , .� �I .� � /� � /� �I .� �I      E  , , -V �� -V Ǳ . Ǳ . �� -V ��      E  , , .� �Y .� �! /� �! /� �Y .� �Y      E  , , -V �I -V � . � . �I -V �I      E  , , -V �	 -V �� . �� . �	 -V �	      E  , , .� �� .� �a /� �a /� �� .� ��      E  , , .� �� .� �� /� �� /� �� .� ��      E  , , .� �� .� �q /� �q /� �� .� ��      E  , , -V �Y -V �! . �! . �Y -V �Y      E  , , .� �� .� Ǳ /� Ǳ /� �� .� ��      E  , , -V �� -V �� . �� . �� -V ��      E  , , .� �i .� �1 /� �1 /� �i .� �i      E  , , -V �� -V �a . �a . �� -V ��      E  , , .� �y .� �A /� �A /� �y .� �y      E  , , -V �� -V �q . �q . �� -V ��      E  , , -V �i -V �1 . �1 . �i -V �i      E  , , .� �� .� �� /� �� /� �� .� ��      E  , , .� �) .� �� /� �� /� �) .� �)      E  , , -V �� -V �� . �� . �� -V ��      E  , , =< W� =< Xj > Xj > W� =< W�      E  , , ;� Y2 ;� Y� <t Y� <t Y2 ;� Y2      E  , , ;� W� ;� Xj <t Xj <t W� ;� W�      E  , , : Y2 : Y� :� Y� :� Y2 : Y2      E  , , : W� : Xj :� Xj :� W� : W�      E  , , A� Y2 A� Y� B� Y� B� Y2 A� Y2      E  , , A� W� A� Xj B� Xj B� W� A� W�      E  , , @\ Y2 @\ Y� A$ Y� A$ Y2 @\ Y2      E  , , @\ W� @\ Xj A$ Xj A$ W� @\ W�      E  , , >� Y2 >� Y� ?� Y� ?� Y2 >� Y2      E  , , >� W� >� Xj ?� Xj ?� W� >� W�      E  , , =< Y2 =< Y� > Y� > Y2 =< Y2      E  , , �\ W� �\ Xj �$ Xj �$ W� �\ W�      E  , , 0� Y2 0� Y� 1� Y� 1� Y2 0� Y2      E  , , � W� � Xj � Xj � W� � W�      E  , , � W� � Xj � Xj � W� � W�      E  , , /, W� /, Xj /� Xj /� W� /, W�      E  , , -� Y2 -� Y� .d Y� .d Y2 -� Y2      E  , , , Y2 , Y� � Y� � Y2 , Y2      E  , , �� Y2 �� Y� �� Y� �� Y2 �� Y2      E  , , l Y2 l Y� 4 Y� 4 Y2 l Y2      E  , , 8� Y2 8� Y� 9T Y� 9T Y2 8� Y2      E  , , \ Y2 \ Y� $ Y� $ Y2 \ Y2      E  , , -� W� -� Xj .d Xj .d W� -� W�      E  , , \ W� \ Xj $ Xj $ W� \ W�      E  , , �� W� �� Xj �� Xj �� W� �� W�      E  , , , Y2 , Y� ,� Y� ,� Y2 , Y2      E  , , � W� � Xj d Xj d W� � W�      E  , ,  Y2  Y� � Y� � Y2  Y2      E  , , 8� W� 8� Xj 9T Xj 9T W� 8� W�      E  , , 6� Y2 6� Y� 7� Y� 7� Y2 6� Y2      E  , , � Y2 � Y� � Y� � Y2 � Y2      E  , , , W� , Xj ,� Xj ,� W� , W�      E  , , *| Y2 *| Y� +D Y� +D Y2 *| Y2      E  , , � W� � Xj � Xj � W� � W�      E  , , � W� � Xj � Xj � W� � W�      E  , , 6� W� 6� Xj 7� Xj 7� W� 6� W�      E  , , � Y2 � Y� � Y� � Y2 � Y2      E  , , � W� � Xj � Xj � W� � W�      E  , , *| W� *| Xj +D Xj +D W� *| W�      E  , , (� Y2 (� Y� )� Y� )� Y2 (� Y2      E  , , 5l Y2 5l Y� 64 Y� 64 Y2 5l Y2      E  , , < Y2 < Y�  Y�  Y2 < Y2      E  , , �, Y2 �, Y� �� Y� �� Y2 �, Y2      E  , , 5l W� 5l Xj 64 Xj 64 W� 5l W�      E  , , < W� < Xj  Xj  W� < W�      E  , , (� W� (� Xj )� Xj )� W� (� W�      E  , , 3� Y2 3� Y� 4� Y� 4� Y2 3� Y2      E  , , �, W� �, Xj �� Xj �� W� �, W�      E  , , '\ Y2 '\ Y� ($ Y� ($ Y2 '\ Y2      E  , , L W� L Xj  Xj  W� L W�      E  , ,  L Y2  L Y�  Y�  Y2  L Y2      E  , , 3� W� 3� Xj 4� Xj 4� W� 3� W�      E  , , 	� Y2 	� Y� 
t Y� 
t Y2 	� Y2      E  , , �� Y2 �� Y� �� Y� �� Y2 �� Y2      E  , , '\ W� '\ Xj ($ Xj ($ W� '\ W�      E  , , %� Y2 %� Y� &� Y� &� Y2 %� Y2      E  , , 2L Y2 2L Y� 3 Y� 3 Y2 2L Y2      E  , ,  L W�  L Xj  Xj  W�  L W�      E  , , 2L W� 2L Xj 3 Xj 3 W� 2L W�      E  , , � Y2 � Y� � Y� � Y2 � Y2      E  , , L Y2 L Y�  Y�  Y2 L Y2      E  , , %� W� %� Xj &� Xj &� W� %� W�      E  , , $< Y2 $< Y� % Y� % Y2 $< Y2      E  , , �� W� �� Xj �� Xj �� W� �� W�      E  , , 	� W� 	� Xj 
t Xj 
t W� 	� W�      E  , , | W� | Xj D Xj D W� | W�      E  , , � W� � Xj � Xj � W� � W�      E  , , l W� l Xj 4 Xj 4 W� l W�      E  , , $< W� $< Xj % Xj % W� $< W�      E  , , �\ Y2 �\ Y� �$ Y� �$ Y2 �\ Y2      E  , ,  W�  Xj � Xj � W�  W�      E  , , "� Y2 "� Y� #t Y� #t Y2 "� Y2      E  , ,  Y2  Y� � Y� � Y2  Y2      E  , , �� Y2 �� Y� �d Y� �d Y2 �� Y2      E  , , �� W� �� Xj �d Xj �d W� �� W�      E  , ,  W�  Xj � Xj � W�  W�      E  , , �| Y2 �| Y� �D Y� �D Y2 �| Y2      E  , , "� W� "� Xj #t Xj #t W� "� W�      E  , , ! Y2 ! Y� !� Y� !� Y2 ! Y2      E  , , �| W� �| Xj �D Xj �D W� �| W�      E  , , | Y2 | Y� D Y� D Y2 | Y2      E  , , , W� , Xj � Xj � W� , W�      E  , , � Y2 � Y� d Y� d Y2 � Y2      E  , , � Y2 � Y� T Y� T Y2 � Y2      E  , , ! W� ! Xj !� Xj !� W� ! W�      E  , , � Y2 � Y�  T Y�  T Y2 � Y2      E  , , � W� � Xj T Xj T W� � W�      E  , , �� W� �� Xj �� Xj �� W� �� W�      E  , , 0� W� 0� Xj 1� Xj 1� W� 0� W�      E  , , l W� l Xj 4 Xj 4 W� l W�      E  , , � Y2 � Y� �� Y� �� Y2 � Y2      E  , , � W� � Xj �� Xj �� W� � W�      E  , , � Y2 � Y� � Y� � Y2 � Y2      E  , , � W� � Xj � Xj � W� � W�      E  , , � W� � Xj  T Xj  T W� � W�      E  , , /, Y2 /, Y� /� Y� /� Y2 /, Y2      E  , , � Y2 � Y� � Y� � Y2 � Y2      E  , , � Y2 � Y� � Y� � Y2 � Y2      E  , , � Y2 � Y� � Y� � Y2 � Y2      E  , , l Y2 l Y� 4 Y� 4 Y2 l Y2      E  , , �� Y2 �� Y� �� Y� �� Y2 �� Y2      E  , ,  @&  @� � @� � @&  @&      E  , , � @& � @� [ @� [ @& � @&      E  , , 
s @& 
s @� ; @� ; @& 
s @&      E  , , � @& � @� 	� @� 	� @& � @&      E  , , 
s QV 
s R ; R ; QV 
s QV      E  , , 
s K 
s K� ; K� ; K 
s K      E  , , � N6 � N� 	� N� 	� N6 � N6      E  , ,  G�  H� � H� � G�  G�      E  , ,  D�  E� � E� � D�  D�      E  , , 
s D� 
s E� ; E� ; D� 
s D�      E  , , � V � V� 	� V� 	� V � V      E  , , � Y& � Y� [ Y� [ Y& � Y&      E  , , � L� � Mn 	� Mn 	� L� � L�      E  , , 
s W� 
s X^ ; X^ ; W� 
s W�      E  , , � Ff � G. [ G. [ Ff � Ff      E  , , 
s Y& 
s Y� ; Y� ; Y& 
s Y&      E  , , 
s Ff 
s G. ; G. ; Ff 
s Ff      E  , ,  V  V� � V� � V  V      E  , , � K � K� 	� K� 	� K � K      E  , , � I� � JN [ JN [ I� � I�      E  , , � W� � X^ [ X^ [ W� � W�      E  , , 
s G� 
s H� ; H� ; G� 
s G�      E  , , 
s A� 
s B~ ; B~ ; A� 
s A�      E  , , � Tv � U> 	� U> 	� Tv � Tv      E  , ,  K  K� � K� � K  K      E  , , 
s N6 
s N� ; N� ; N6 
s N6      E  , , � O� � P� [ P� [ O� � O�      E  , , � D� � E� [ E� [ D� � D�      E  , , � I� � JN 	� JN 	� I� � I�      E  , , � O� � P� 	� P� 	� O� � O�      E  , , � A� � B~ 	� B~ 	� A� � A�      E  , , � V � V� [ V� [ V � V      E  , ,  CF  D � D � CF  CF      E  , ,  I�  JN � JN � I�  I�      E  , , � G� � H� 	� H� 	� G� � G�      E  , , � Tv � U> [ U> [ Tv � Tv      E  , ,  W�  X^ � X^ � W�  W�      E  , , 
s Tv 
s U> ; U> ; Tv 
s Tv      E  , ,  Tv  U> � U> � Tv  Tv      E  , , 
s I� 
s JN ; JN ; I� 
s I�      E  , , � R� � S� 	� S� 	� R� � R�      E  , , � Ff � G. 	� G. 	� Ff � Ff      E  , ,  N6  N� � N� � N6  N6      E  , , � CF � D [ D [ CF � CF      E  , , 
s V 
s V� ; V� ; V 
s V      E  , , 
s R� 
s S� ; S� ; R� 
s R�      E  , ,  Y&  Y� � Y� � Y&  Y&      E  , , 
s L� 
s Mn ; Mn ; L� 
s L�      E  , , � Y& � Y� 	� Y� 	� Y& � Y&      E  , , � R� � S� [ S� [ R� � R�      E  , ,  Ff  G. � G. � Ff  Ff      E  , , � D� � E� 	� E� 	� D� � D�      E  , , 
s O� 
s P� ; P� ; O� 
s O�      E  , , 
s CF 
s D ; D ; CF 
s CF      E  , , � A� � B~ [ B~ [ A� � A�      E  , , � G� � H� [ H� [ G� � G�      E  , ,  QV  R � R � QV  QV      E  , , � CF � D 	� D 	� CF � CF      E  , , � QV � R [ R [ QV � QV      E  , ,  O�  P� � P� � O�  O�      E  , ,  A�  B~ � B~ � A�  A�      E  , , � K � K� [ K� [ K � K      E  , ,  L�  Mn � Mn � L�  L�      E  , , � L� � Mn [ Mn [ L� � L�      E  , ,  R�  S� � S� � R�  R�      E  , , � QV � R 	� R 	� QV � QV      E  , , � W� � X^ 	� X^ 	� W� � W�      E  , , � N6 � N� [ N� [ N6 � N6      E  , , 
s 6� 
s 7� ; 7� ; 6� 
s 6�      E  , , � 6� � 7� 	� 7� 	� 6� � 6�      E  , ,  %�  &^ � &^ � %�  %�      E  , , 
s = 
s =� ; =� ; = 
s =      E  , ,  +�  ,� � ,� � +�  +�      E  , , � 56 � 5� [ 5� [ 56 � 56      E  , , � 3� � 4n 	� 4n 	� 3� � 3�      E  , ,  >�  ?^ � ?^ � >�  >�      E  , , � 0� � 1N [ 1N [ 0� � 0�      E  , , 
s ;v 
s <> ; <> ; ;v 
s ;v      E  , , � 9� � :� 	� :� 	� 9� � 9�      E  , , 
s %� 
s &^ ; &^ ; %� 
s %�      E  , , � 56 � 5� 	� 5� 	� 56 � 56      E  , , � (� � )~ [ )~ [ (� � (�      E  , , � '& � '� [ '� [ '& � '&      E  , , � -f � .. 	� .. 	� -f � -f      E  , , � *F � + 	� + 	� *F � *F      E  , , 
s 9� 
s :� ; :� ; 9� 
s 9�      E  , , � 0� � 1N 	� 1N 	� 0� � 0�      E  , , 
s .� 
s /� ; /� ; .� 
s .�      E  , , � ;v � <> [ <> [ ;v � ;v      E  , , 
s 8V 
s 9 ; 9 ; 8V 
s 8V      E  , ,  9�  :� � :� � 9�  9�      E  , , � 8V � 9 	� 9 	� 8V � 8V      E  , , 
s 3� 
s 4n ; 4n ; 3� 
s 3�      E  , , � 9� � :� [ :� [ 9� � 9�      E  , ,  0�  1N � 1N � 0�  0�      E  , , � .� � /� [ /� [ .� � .�      E  , , 
s 56 
s 5� ; 5� ; 56 
s 56      E  , , � >� � ?^ [ ?^ [ >� � >�      E  , ,  6�  7� � 7� � 6�  6�      E  , , � *F � + [ + [ *F � *F      E  , , 
s *F 
s + ; + ; *F 
s *F      E  , ,  -f  .. � .. � -f  -f      E  , ,  3�  4n � 4n � 3�  3�      E  , , � = � =� [ =� [ = � =      E  , , 
s (� 
s )~ ; )~ ; (� 
s (�      E  , ,  =  =� � =� � =  =      E  , ,  *F  + � + � *F  *F      E  , , � 2 � 2� 	� 2� 	� 2 � 2      E  , ,  56  5� � 5� � 56  56      E  , ,  .�  /� � /� � .�  .�      E  , , � 8V � 9 [ 9 [ 8V � 8V      E  , , � +� � ,� [ ,� [ +� � +�      E  , ,  (�  )~ � )~ � (�  (�      E  , , � -f � .. [ .. [ -f � -f      E  , , 
s -f 
s .. ; .. ; -f 
s -f      E  , , � 2 � 2� [ 2� [ 2 � 2      E  , , � +� � ,� 	� ,� 	� +� � +�      E  , ,  8V  9 � 9 � 8V  8V      E  , , � '& � '� 	� '� 	� '& � '&      E  , , 
s 0� 
s 1N ; 1N ; 0� 
s 0�      E  , , � >� � ?^ 	� ?^ 	� >� � >�      E  , , 
s 2 
s 2� ; 2� ; 2 
s 2      E  , , 
s +� 
s ,� ; ,� ; +� 
s +�      E  , , � 6� � 7� [ 7� [ 6� � 6�      E  , , 
s '& 
s '� ; '� ; '& 
s '&      E  , ,  ;v  <> � <> � ;v  ;v      E  , , � (� � )~ 	� )~ 	� (� � (�      E  , , � = � =� 	� =� 	� = � =      E  , , � 3� � 4n [ 4n [ 3� � 3�      E  , , � %� � &^ [ &^ [ %� � %�      E  , , � ;v � <> 	� <> 	� ;v � ;v      E  , , � %� � &^ 	� &^ 	� %� � %�      E  , ,  '&  '� � '� � '&  '&      E  , , 
s >� 
s ?^ ; ?^ ; >� 
s >�      E  , ,  2  2� � 2� � 2  2      E  , , � .� � /� 	� /� 	� .� � .�      E  , , � 	v � 
> [ 
> [ 	v � 	v      E  , ,  	v  
> � 
> � 	v  	v      E  , , � 	v � 
> 	� 
> 	� 	v � 	v      E  , , 
s 	v 
s 
> ; 
> ; 	v 
s 	v      E  , , 
s � 
s N ; N ; � 
s �      E  , ,  �  ~ � ~ � �  �      E  , , � V �   [   [ V � V      E  , , � � � � 	� � 	� � � �      E  , , � "v � #> [ #> [ "v � "v      E  , , 
s � 
s ^ ; ^ ; � 
s �      E  , , � � � n 	� n 	� � � �      E  , , � � � � 	� � 	� � � �      E  , , �  � � [ � [  �       E  , , � F �  	�  	� F � F      E  , , �  � � [ � [  �       E  , , 
s  � 
s !� ; !� ;  � 
s  �      E  , , 
s & 
s � ; � ; & 
s &      E  , , � � � N 	� N 	� � � �      E  , , 
s V 
s   ;   ; V 
s V      E  , ,  �  N � N � �  �      E  , , 
s � 
s � ; � ; � 
s �      E  , , � � � n [ n [ � � �      E  , , � $ � $� [ $� [ $ � $      E  , , � $ � $� 	� $� 	� $ � $      E  , ,  &  � � � � &  &      E  , ,  f  . � . � f  f      E  , , 
s 6 
s � ; � ; 6 
s 6      E  , , � � � � [ � [ � � �      E  , , 
s f 
s . ; . ; f 
s f      E  , ,  F   �  � F  F      E  , ,  �  n � n � �  �      E  , , � f � . [ . [ f � f      E  , ,   �  !� � !� �  �   �      E  , , � V �   	�   	� V � V      E  , , � f � . 	� . 	� f � f      E  , ,  �  � � � � �  �      E  , , � F �  [  [ F � F      E  , , � 6 � � 	� � 	� 6 � 6      E  , , 
s  
s � ; � ;  
s       E  , , 
s "v 
s #> ; #> ; "v 
s "v      E  , , 
s  
s � ; � ;  
s       E  , ,  "v  #> � #> � "v  "v      E  , ,  �  � � � � �  �      E  , , � "v � #> 	� #> 	� "v � "v      E  , , � � � ^ [ ^ [ � � �      E  , , � � � � [ � [ � � �      E  , ,  $  $� � $� � $  $      E  , , � � � ^ 	� ^ 	� � � �      E  , , 
s F 
s  ;  ; F 
s F      E  , , � & � � 	� � 	� & � &      E  , , 
s $ 
s $� ; $� ; $ 
s $      E  , ,  6  � � � � 6  6      E  , , �  � � !� [ !� [  � �  �      E  , , � � � N [ N [ � � �      E  , , �  � � !� 	� !� 	�  � �  �      E  , , 
s � 
s ~ ; ~ ; � 
s �      E  , , � & � � [ � [ & � &      E  , , � � � ~ 	� ~ 	� � � �      E  , ,    � � � �         E  , , 
s � 
s � ; � ; � 
s �      E  , ,  �  � � � � �  �      E  , ,  V    �   � V  V      E  , ,    � � � �         E  , , 
s � 
s � ; � ; � 
s �      E  , , � � � � [ � [ � � �      E  , , � � � ~ [ ~ [ � � �      E  , , �  � � 	� � 	�  �       E  , , � 6 � � [ � [ 6 � 6      E  , , �  � � 	� � 	�  �       E  , , 
s � 
s n ; n ; � 
s �      E  , , � � � � 	� � 	� � � �      E  , ,  �  ^ � ^ � �  �      E  , , �  �� �  �~ 	�  �~ 	�  �� �  ��      E  , , 
s  �F 
s  � ;  � ;  �F 
s  �F      E  , ,   �f   �. �  �. �  �f   �f      E  , ,      � �  � �           E  , , �  �� �  �N 	�  �N 	�  �� �  ��      E  , , �  � �  �� 	�  �� 	�  � �  �      E  , , 
s   
s  � ;  � ;   
s        E  , ,  6  � � � � 6  6      E  , ,   ��   �~ �  �~ �  ��   ��      E  , , �  �F �  � 	�  � 	�  �F �  �F      E  , , �  � �  �^ [  �^ [  � �  �      E  , , � � � n [ n [ � � �      E  , , �  �F �  � [  � [  �F �  �F      E  , , �  �& �  �� [  �� [  �& �  �&      E  , , 
s � 
s � ; � ; � 
s �      E  , ,   ��   �� �  �� �  ��   ��      E  , , � � � n 	� n 	� � � �      E  , , �  �v �  �> 	�  �> 	�  �v �  �v      E  , , �  �v �  �> [  �> [  �v �  �v      E  , , �  � �  �� [  �� [  � �  �      E  , , 
s  �� 
s  �� ;  �� ;  �� 
s  ��      E  , ,   �   �� �  �� �  �   �      E  , ,  �  � � � � �  �      E  , , � 6 � � [ � [ 6 � 6      E  , , 
s V 
s  ;  ; V 
s V      E  , , � � � � 	� � 	� � � �      E  , ,  V   �  � V  V      E  , , �  �f �  �. 	�  �. 	�  �f �  �f      E  , , �  �� �  �� 	�  �� 	�  �� �  ��      E  , ,  �  � � � � �  �      E  , , �  �� �  �� [  �� [  �� �  ��      E  , , � V �  	�  	� V � V      E  , , �  �� �  � 	�  � 	�  �� �  ��      E  , , 
s  �� 
s  �~ ;  �~ ;  �� 
s  ��      E  , , �   �  � [  � [   �        E  , ,   �&   �� �  �� �  �&   �&      E  , ,   ��   � �  � �  ��   ��      E  , , �  �& �  �� 	�  �� 	�  �& �  �&      E  , , 
s � 
s � ; � ; � 
s �      E  , , 
s  �f 
s  �. ;  �. ;  �f 
s  �f      E  , ,   �F   � �  � �  �F   �F      E  , , 
s  �& 
s  �� ;  �� ;  �& 
s  �&      E  , , 
s  �� 
s  � ;  � ;  �� 
s  ��      E  , , �  �� �  �� 	�  �� 	�  �� �  ��      E  , ,   ��   �� �  �� �  ��   ��      E  , , �  �� �  �~ [  �~ [  �� �  ��      E  , , �  �f �  �. [  �. [  �f �  �f      E  , , �   �  � 	�  � 	�   �        E  , ,   �v   �> �  �> �  �v   �v      E  , , �  � �  �^ 	�  �^ 	�  � �  �      E  , , � V �  [  [ V � V      E  , , 
s  � 
s  �� ;  �� ;  � 
s  �      E  , , 
s � 
s n ; n ; � 
s �      E  , , �  �� �  �N [  �N [  �� �  ��      E  , , �  �� �  �� [  �� [  �� �  ��      E  , ,   ��   �N �  �N �  ��   ��      E  , , 
s  �v 
s  �> ;  �> ;  �v 
s  �v      E  , , � � � � [ � [ � � �      E  , , 
s  �� 
s  �N ;  �N ;  �� 
s  ��      E  , , 
s  �� 
s  �� ;  �� ;  �� 
s  ��      E  , , � � � � [ � [ � � �      E  , ,   �   �^ �  �^ �  �   �      E  , , 
s 6 
s � ; � ; 6 
s 6      E  , , �  �� �  � [  � [  �� �  ��      E  , , � � � � 	� � 	� � � �      E  , , � 6 � � 	� � 	� 6 � 6      E  , , 
s  � 
s  �^ ;  �^ ;  � 
s  �      E  , ,  �  n � n � �  �      G   ,  ��  ��  �� ��  �� ��  ��  ��  ��  ��      G   , �  �� � �� � �� �  �� �  ��      F   ,  �� �B  �� �� I� �� I� �B  �� �B      F   , K� |@ K� }� T+ }� T+ |@ K� |@      F   ,  ��  ��  �� �B �L �B �L  ��  ��  ��      F   ,  �� �B  �� ��  �� ��  �� �B  �� �B      F   , �9 �B �9 �� �L �� �L �B �9 �B      F   , �  �� � �� � �� �  �� �  ��      G   , �  �� � �� � �� �  �� �  ��      G   , �� �� �� �� � �� � �� �� ��      G   , �� �� �� �� �� �� �� �� �� ��      G   , � �� � �� �I �� �I �� � ��      G   , �U �� �U �� �� �� �� �� �U ��      G   , �� �� �� �� �� �� �� �� �� ��      G   , �� �� �� �� �� �� �� �� �� ��      G   , �� �� �� �� �) �� �) �� �� ��      G   , v5 �� v5 �� wa �� wa �� v5 ��      G   , km �� km �� l� �� l� �� km ��      G   , `� �� `� �� a� �� a� �� `� ��      G   , U� �� U� �� W	 �� W	 �� U� ��      G   , K �� K �� LA �� LA �� K ��      G   , @M �� @M �� Ay �� Ay �� @M ��      G   , 5� �� 5� �� 6� �� 6� �� 5� ��      G   , *� �� *� �� +� �� +� �� *� ��      G   , � �� � �� !! �� !! �� � ��      G   , - �� - �� Y �� Y �� - ��      G   , 
e �� 
e �� � �� � �� 
e ��      G   , �� �� �� ��  � ��  � �� �� ��      G   , HU �� HU �� I� �� I� �� HU ��      G   , =� �� =� �� >� �� >� �� =� ��      G   , 2� �� 2� �� 3� �� 3� �� 2� ��      G   , '� �� '� �� )) �� )) �� '� ��      G   , 5 �� 5 �� a �� a �� 5 ��      G   , m �� m �� � �� � �� m ��      G   , � �� � �� � �� � �� � ��      G   ,  �� ��  �� ��  �	 ��  �	 ��  �� ��      G   , �� �� �� �� �� �� �� �� �� ��      G   , �� �� �� �� �� �� �� �� �� ��      G   , � �� � �� �1 �� �1 �� � ��      G   , ~= �� ~= �� i �� i �� ~= ��      G   , su �� su �� t� �� t� �� su ��      G   , h� �� h� �� i� �� i� �� h� ��      G   , ]� �� ]� �� _ �� _ �� ]� ��      G   , S �� S �� TI �� TI �� S ��      G   , �� �� �� �� � �� � �� �� ��      G   , � �� � �� �9 �� �9 �� � ��      G   , �E �� �E �� �q �� �q �� �E ��      G   , �} �� �} �� թ �� թ �� �} ��      G   ,  ��  ��  �� ��  �� ��  ��  ��  ��  ��      G   , ɵ �� ɵ �� �� �� �� �� ɵ ��      G   , �� �� �� �� � �� � �� �� ��      G   , �% �� �% �� �Q �� �Q �� �% ��      G   , �] �� �] �� �� �� �� �� �] ��      G        A        � Ѭ VGND      G    �{ �� clk       G    �C �� ena       G    �� �� 
rst_n       G    �� �� ui_in[0]      G    �# �� ui_in[1]      G    �[ �� ui_in[2]      G    �� �� ui_in[3]      G    v� �� ui_in[4]      G    l �� ui_in[5]      G    a; �� ui_in[6]      G    Vs �� ui_in[7]      G    K� �� uio_in[0]       G    @� �� uio_in[1]       G    6 �� uio_in[2]       G    +S �� uio_in[3]       G     � �� uio_in[4]       G    � �� uio_in[5]       G    
� �� uio_in[6]       G     3 �� uio_in[7]       G    H� �� uio_oe[0]       G    ># �� uio_oe[1]       G    3[ �� uio_oe[2]       G    (� �� uio_oe[3]       G    � �� uio_oe[4]       G     �� uio_oe[5]       G    ; �� uio_oe[6]       G     �s �� uio_oe[7]       G    �+ �� uio_out[0]      G    �c �� uio_out[1]      G    �� �� uio_out[2]      G    ~� �� uio_out[3]      G    t �� uio_out[4]      G    iC �� uio_out[5]      G    ^{ �� uio_out[6]      G    S� �� uio_out[7]      G    �k �� uo_out[0]       G    � �� uo_out[1]       G    �� �� uo_out[2]       G    � �� uo_out[3]       G    �K �� uo_out[4]       G    �� �� uo_out[5]       G    �� �� uo_out[6]       G    �� �� uo_out[7]       G        A         �Y � VPWR      