VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_wulf_8bit_vco
  CLASS BLOCK ;
  FOREIGN tt_um_wulf_8bit_vco ;
  ORIGIN -43.263 -60.898 ;
  SIZE 157.320 BY 111.520 ;
END tt_um_wulf_8bit_vco
END LIBRARY

