VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_wulf_8bit_vco
  CLASS BLOCK ;
  FOREIGN tt_um_wulf_8bit_vco ;
  ORIGIN 0.000 0.000 ;
  SIZE 157.320 BY 111.520 ;
  PIN VGND
    ANTENNADIFFAREA 5.390300 ;
    PORT
      LAYER li1 ;
        RECT 85.455 106.355 102.475 106.525 ;
        RECT 85.990 105.875 86.160 106.355 ;
        RECT 86.830 105.875 87.000 106.355 ;
        RECT 87.670 105.875 87.840 106.355 ;
        RECT 88.510 105.875 88.680 106.355 ;
        RECT 89.350 105.875 89.520 106.355 ;
        RECT 90.190 105.875 90.360 106.355 ;
        RECT 91.030 105.875 91.200 106.355 ;
        RECT 91.870 105.875 92.040 106.355 ;
        RECT 92.710 105.875 92.880 106.355 ;
        RECT 93.550 105.875 93.720 106.355 ;
        RECT 94.390 105.875 94.560 106.355 ;
        RECT 95.230 105.535 95.400 106.355 ;
        RECT 96.050 105.555 96.380 106.355 ;
        RECT 96.890 105.875 97.220 106.355 ;
        RECT 97.730 105.875 98.060 106.355 ;
        RECT 98.570 105.875 98.900 106.355 ;
        RECT 99.410 105.875 99.740 106.355 ;
        RECT 100.250 105.875 100.580 106.355 ;
        RECT 101.620 105.975 101.950 106.355 ;
        RECT 11.625 102.050 12.315 102.220 ;
        RECT 129.710 101.990 131.890 102.340 ;
        RECT 56.855 100.150 57.545 100.320 ;
        RECT 111.545 88.515 111.715 89.205 ;
        RECT 6.130 47.990 6.300 48.680 ;
        RECT 105.530 16.485 106.220 16.655 ;
        RECT 65.315 6.890 66.005 7.060 ;
        RECT 12.180 5.735 12.350 6.425 ;
      LAYER mcon ;
        RECT 85.600 106.355 85.770 106.525 ;
        RECT 86.060 106.355 86.230 106.525 ;
        RECT 86.520 106.355 86.690 106.525 ;
        RECT 86.980 106.355 87.150 106.525 ;
        RECT 87.440 106.355 87.610 106.525 ;
        RECT 87.900 106.355 88.070 106.525 ;
        RECT 88.360 106.355 88.530 106.525 ;
        RECT 88.820 106.355 88.990 106.525 ;
        RECT 89.280 106.355 89.450 106.525 ;
        RECT 89.740 106.355 89.910 106.525 ;
        RECT 90.200 106.355 90.370 106.525 ;
        RECT 90.660 106.355 90.830 106.525 ;
        RECT 91.120 106.355 91.290 106.525 ;
        RECT 91.580 106.355 91.750 106.525 ;
        RECT 92.040 106.355 92.210 106.525 ;
        RECT 92.500 106.355 92.670 106.525 ;
        RECT 92.960 106.355 93.130 106.525 ;
        RECT 93.420 106.355 93.590 106.525 ;
        RECT 93.880 106.355 94.050 106.525 ;
        RECT 94.340 106.355 94.510 106.525 ;
        RECT 94.800 106.355 94.970 106.525 ;
        RECT 95.260 106.355 95.430 106.525 ;
        RECT 95.720 106.355 95.890 106.525 ;
        RECT 96.180 106.355 96.350 106.525 ;
        RECT 96.640 106.355 96.810 106.525 ;
        RECT 97.100 106.355 97.270 106.525 ;
        RECT 97.560 106.355 97.730 106.525 ;
        RECT 98.020 106.355 98.190 106.525 ;
        RECT 98.480 106.355 98.650 106.525 ;
        RECT 98.940 106.355 99.110 106.525 ;
        RECT 99.400 106.355 99.570 106.525 ;
        RECT 99.860 106.355 100.030 106.525 ;
        RECT 100.320 106.355 100.490 106.525 ;
        RECT 100.780 106.355 100.950 106.525 ;
        RECT 101.240 106.355 101.410 106.525 ;
        RECT 101.700 106.355 101.870 106.525 ;
        RECT 102.160 106.355 102.330 106.525 ;
        RECT 11.705 102.050 11.875 102.220 ;
        RECT 12.065 102.050 12.235 102.220 ;
        RECT 129.820 102.080 129.990 102.250 ;
        RECT 130.180 102.080 130.350 102.250 ;
        RECT 130.540 102.080 130.710 102.250 ;
        RECT 130.900 102.080 131.070 102.250 ;
        RECT 131.260 102.080 131.430 102.250 ;
        RECT 131.620 102.080 131.790 102.250 ;
        RECT 56.935 100.150 57.105 100.320 ;
        RECT 57.295 100.150 57.465 100.320 ;
        RECT 111.545 88.955 111.715 89.125 ;
        RECT 111.545 88.595 111.715 88.765 ;
        RECT 6.130 48.430 6.300 48.600 ;
        RECT 6.130 48.070 6.300 48.240 ;
        RECT 105.610 16.485 105.780 16.655 ;
        RECT 105.970 16.485 106.140 16.655 ;
        RECT 65.395 6.890 65.565 7.060 ;
        RECT 65.755 6.890 65.925 7.060 ;
        RECT 12.180 6.175 12.350 6.345 ;
        RECT 12.180 5.815 12.350 5.985 ;
      LAYER met1 ;
        RECT 21.435 108.930 21.805 109.650 ;
        RECT 24.195 108.930 24.565 109.650 ;
        RECT 26.955 108.930 27.325 109.650 ;
        RECT 29.715 108.930 30.085 109.650 ;
        RECT 32.475 108.930 32.845 109.650 ;
        RECT 35.235 108.930 35.605 109.650 ;
        RECT 37.995 108.930 38.365 109.650 ;
        RECT 40.755 108.930 41.125 109.650 ;
        RECT 43.515 108.930 43.885 109.650 ;
        RECT 46.275 108.930 46.645 109.650 ;
        RECT 49.035 108.930 49.405 109.650 ;
        RECT 51.795 108.930 52.165 109.650 ;
        RECT 54.555 108.930 54.925 109.650 ;
        RECT 57.315 108.930 57.685 109.650 ;
        RECT 60.075 108.930 60.445 109.650 ;
        RECT 62.835 108.930 63.205 109.650 ;
        RECT 65.595 108.930 65.965 109.650 ;
        RECT 68.355 108.930 68.725 109.650 ;
        RECT 71.115 108.930 71.485 109.650 ;
        RECT 73.875 108.930 74.245 109.650 ;
        RECT 76.635 108.930 77.005 109.650 ;
        RECT 79.395 108.930 79.765 109.650 ;
        RECT 82.155 108.930 82.525 109.650 ;
        RECT 85.455 106.200 102.475 106.680 ;
        RECT 13.245 102.755 13.505 103.015 ;
        RECT 13.645 102.755 13.905 103.015 ;
        RECT 14.045 102.755 14.305 103.015 ;
        RECT 14.445 102.755 14.705 103.015 ;
        RECT 14.845 102.755 15.105 103.015 ;
        RECT 15.245 102.755 15.505 103.015 ;
        RECT 15.645 102.755 15.905 103.015 ;
        RECT 16.045 102.755 16.305 103.015 ;
        RECT 16.445 102.755 16.705 103.015 ;
        RECT 16.845 102.755 17.105 103.015 ;
        RECT 17.245 102.755 17.505 103.015 ;
        RECT 17.645 102.755 17.905 103.015 ;
        RECT 13.245 102.355 13.505 102.615 ;
        RECT 13.645 102.355 13.905 102.615 ;
        RECT 14.045 102.355 14.305 102.615 ;
        RECT 14.445 102.355 14.705 102.615 ;
        RECT 14.845 102.355 15.105 102.615 ;
        RECT 15.245 102.355 15.505 102.615 ;
        RECT 15.645 102.355 15.905 102.615 ;
        RECT 16.045 102.355 16.305 102.615 ;
        RECT 16.445 102.355 16.705 102.615 ;
        RECT 16.845 102.355 17.105 102.615 ;
        RECT 17.245 102.355 17.505 102.615 ;
        RECT 17.645 102.355 17.905 102.615 ;
        RECT 11.630 102.020 12.310 102.340 ;
        RECT 129.745 102.005 131.865 102.325 ;
        RECT 58.510 100.905 58.770 101.165 ;
        RECT 58.910 100.905 59.170 101.165 ;
        RECT 59.310 100.905 59.570 101.165 ;
        RECT 59.710 100.905 59.970 101.165 ;
        RECT 60.110 100.905 60.370 101.165 ;
        RECT 60.510 100.905 60.770 101.165 ;
        RECT 60.910 100.905 61.170 101.165 ;
        RECT 61.310 100.905 61.570 101.165 ;
        RECT 61.710 100.905 61.970 101.165 ;
        RECT 62.110 100.905 62.370 101.165 ;
        RECT 62.510 100.905 62.770 101.165 ;
        RECT 62.910 100.905 63.170 101.165 ;
        RECT 58.510 100.505 58.770 100.765 ;
        RECT 58.910 100.505 59.170 100.765 ;
        RECT 59.310 100.505 59.570 100.765 ;
        RECT 59.710 100.505 59.970 100.765 ;
        RECT 60.110 100.505 60.370 100.765 ;
        RECT 60.510 100.505 60.770 100.765 ;
        RECT 60.910 100.505 61.170 100.765 ;
        RECT 61.310 100.505 61.570 100.765 ;
        RECT 61.710 100.505 61.970 100.765 ;
        RECT 62.110 100.505 62.370 100.765 ;
        RECT 62.510 100.505 62.770 100.765 ;
        RECT 62.910 100.505 63.170 100.765 ;
        RECT 56.860 100.120 57.540 100.440 ;
        RECT 111.515 88.520 111.835 89.200 ;
        RECT 111.845 87.290 112.105 87.550 ;
        RECT 112.245 87.290 112.505 87.550 ;
        RECT 111.845 86.890 112.105 87.150 ;
        RECT 112.245 86.890 112.505 87.150 ;
        RECT 111.845 86.490 112.105 86.750 ;
        RECT 112.245 86.490 112.505 86.750 ;
        RECT 111.845 86.090 112.105 86.350 ;
        RECT 112.245 86.090 112.505 86.350 ;
        RECT 111.845 85.690 112.105 85.950 ;
        RECT 112.245 85.690 112.505 85.950 ;
        RECT 111.845 85.290 112.105 85.550 ;
        RECT 112.245 85.290 112.505 85.550 ;
        RECT 111.845 84.890 112.105 85.150 ;
        RECT 112.245 84.890 112.505 85.150 ;
        RECT 111.845 84.490 112.105 84.750 ;
        RECT 112.245 84.490 112.505 84.750 ;
        RECT 111.845 84.090 112.105 84.350 ;
        RECT 112.245 84.090 112.505 84.350 ;
        RECT 111.845 83.690 112.105 83.950 ;
        RECT 112.245 83.690 112.505 83.950 ;
        RECT 111.845 83.290 112.105 83.550 ;
        RECT 112.245 83.290 112.505 83.550 ;
        RECT 111.845 82.890 112.105 83.150 ;
        RECT 112.245 82.890 112.505 83.150 ;
        RECT 5.305 54.020 5.565 54.280 ;
        RECT 5.705 54.020 5.965 54.280 ;
        RECT 5.305 53.620 5.565 53.880 ;
        RECT 5.705 53.620 5.965 53.880 ;
        RECT 5.305 53.220 5.565 53.480 ;
        RECT 5.705 53.220 5.965 53.480 ;
        RECT 5.305 52.820 5.565 53.080 ;
        RECT 5.705 52.820 5.965 53.080 ;
        RECT 5.305 52.420 5.565 52.680 ;
        RECT 5.705 52.420 5.965 52.680 ;
        RECT 5.305 52.020 5.565 52.280 ;
        RECT 5.705 52.020 5.965 52.280 ;
        RECT 5.305 51.620 5.565 51.880 ;
        RECT 5.705 51.620 5.965 51.880 ;
        RECT 5.305 51.220 5.565 51.480 ;
        RECT 5.705 51.220 5.965 51.480 ;
        RECT 5.305 50.820 5.565 51.080 ;
        RECT 5.705 50.820 5.965 51.080 ;
        RECT 5.305 50.420 5.565 50.680 ;
        RECT 5.705 50.420 5.965 50.680 ;
        RECT 5.305 50.020 5.565 50.280 ;
        RECT 5.705 50.020 5.965 50.280 ;
        RECT 5.305 49.620 5.565 49.880 ;
        RECT 5.705 49.620 5.965 49.880 ;
        RECT 6.010 47.995 6.330 48.675 ;
        RECT 105.535 16.365 106.215 16.685 ;
        RECT 99.930 16.075 100.190 16.335 ;
        RECT 100.330 16.075 100.590 16.335 ;
        RECT 100.730 16.075 100.990 16.335 ;
        RECT 101.130 16.075 101.390 16.335 ;
        RECT 101.530 16.075 101.790 16.335 ;
        RECT 101.930 16.075 102.190 16.335 ;
        RECT 102.330 16.075 102.590 16.335 ;
        RECT 102.730 16.075 102.990 16.335 ;
        RECT 103.130 16.075 103.390 16.335 ;
        RECT 103.530 16.075 103.790 16.335 ;
        RECT 103.930 16.075 104.190 16.335 ;
        RECT 104.330 16.075 104.590 16.335 ;
        RECT 99.930 15.675 100.190 15.935 ;
        RECT 100.330 15.675 100.590 15.935 ;
        RECT 100.730 15.675 100.990 15.935 ;
        RECT 101.130 15.675 101.390 15.935 ;
        RECT 101.530 15.675 101.790 15.935 ;
        RECT 101.930 15.675 102.190 15.935 ;
        RECT 102.330 15.675 102.590 15.935 ;
        RECT 102.730 15.675 102.990 15.935 ;
        RECT 103.130 15.675 103.390 15.935 ;
        RECT 103.530 15.675 103.790 15.935 ;
        RECT 103.930 15.675 104.190 15.935 ;
        RECT 104.330 15.675 104.590 15.935 ;
        RECT 11.280 11.820 11.540 12.080 ;
        RECT 11.680 11.820 11.940 12.080 ;
        RECT 11.280 11.420 11.540 11.680 ;
        RECT 11.680 11.420 11.940 11.680 ;
        RECT 11.280 11.020 11.540 11.280 ;
        RECT 11.680 11.020 11.940 11.280 ;
        RECT 11.280 10.620 11.540 10.880 ;
        RECT 11.680 10.620 11.940 10.880 ;
        RECT 11.280 10.220 11.540 10.480 ;
        RECT 11.680 10.220 11.940 10.480 ;
        RECT 11.280 9.820 11.540 10.080 ;
        RECT 11.680 9.820 11.940 10.080 ;
        RECT 11.280 9.420 11.540 9.680 ;
        RECT 11.680 9.420 11.940 9.680 ;
        RECT 11.280 9.020 11.540 9.280 ;
        RECT 11.680 9.020 11.940 9.280 ;
        RECT 11.280 8.620 11.540 8.880 ;
        RECT 11.680 8.620 11.940 8.880 ;
        RECT 11.280 8.220 11.540 8.480 ;
        RECT 11.680 8.220 11.940 8.480 ;
        RECT 11.280 7.820 11.540 8.080 ;
        RECT 11.680 7.820 11.940 8.080 ;
        RECT 11.280 7.420 11.540 7.680 ;
        RECT 11.680 7.420 11.940 7.680 ;
        RECT 65.320 6.770 66.000 7.090 ;
        RECT 59.720 6.505 59.980 6.765 ;
        RECT 60.120 6.505 60.380 6.765 ;
        RECT 60.520 6.505 60.780 6.765 ;
        RECT 60.920 6.505 61.180 6.765 ;
        RECT 61.320 6.505 61.580 6.765 ;
        RECT 61.720 6.505 61.980 6.765 ;
        RECT 62.120 6.505 62.380 6.765 ;
        RECT 62.520 6.505 62.780 6.765 ;
        RECT 62.920 6.505 63.180 6.765 ;
        RECT 63.320 6.505 63.580 6.765 ;
        RECT 63.720 6.505 63.980 6.765 ;
        RECT 64.120 6.505 64.380 6.765 ;
        RECT 12.060 5.740 12.380 6.420 ;
        RECT 59.720 6.105 59.980 6.365 ;
        RECT 60.120 6.105 60.380 6.365 ;
        RECT 60.520 6.105 60.780 6.365 ;
        RECT 60.920 6.105 61.180 6.365 ;
        RECT 61.320 6.105 61.580 6.365 ;
        RECT 61.720 6.105 61.980 6.365 ;
        RECT 62.120 6.105 62.380 6.365 ;
        RECT 62.520 6.105 62.780 6.365 ;
        RECT 62.920 6.105 63.180 6.365 ;
        RECT 63.320 6.105 63.580 6.365 ;
        RECT 63.720 6.105 63.980 6.365 ;
        RECT 64.120 6.105 64.380 6.365 ;
      LAYER via ;
        RECT 21.490 109.335 21.750 109.595 ;
        RECT 21.490 108.985 21.750 109.245 ;
        RECT 24.250 109.335 24.510 109.595 ;
        RECT 24.250 108.985 24.510 109.245 ;
        RECT 27.010 109.335 27.270 109.595 ;
        RECT 27.010 108.985 27.270 109.245 ;
        RECT 29.770 109.335 30.030 109.595 ;
        RECT 29.770 108.985 30.030 109.245 ;
        RECT 32.530 109.335 32.790 109.595 ;
        RECT 32.530 108.985 32.790 109.245 ;
        RECT 35.290 109.335 35.550 109.595 ;
        RECT 35.290 108.985 35.550 109.245 ;
        RECT 38.050 109.335 38.310 109.595 ;
        RECT 38.050 108.985 38.310 109.245 ;
        RECT 40.810 109.335 41.070 109.595 ;
        RECT 40.810 108.985 41.070 109.245 ;
        RECT 43.570 109.335 43.830 109.595 ;
        RECT 43.570 108.985 43.830 109.245 ;
        RECT 46.330 109.335 46.590 109.595 ;
        RECT 46.330 108.985 46.590 109.245 ;
        RECT 49.090 109.335 49.350 109.595 ;
        RECT 49.090 108.985 49.350 109.245 ;
        RECT 51.850 109.335 52.110 109.595 ;
        RECT 51.850 108.985 52.110 109.245 ;
        RECT 54.610 109.335 54.870 109.595 ;
        RECT 54.610 108.985 54.870 109.245 ;
        RECT 57.370 109.335 57.630 109.595 ;
        RECT 57.370 108.985 57.630 109.245 ;
        RECT 60.130 109.335 60.390 109.595 ;
        RECT 60.130 108.985 60.390 109.245 ;
        RECT 62.890 109.335 63.150 109.595 ;
        RECT 62.890 108.985 63.150 109.245 ;
        RECT 65.650 109.335 65.910 109.595 ;
        RECT 65.650 108.985 65.910 109.245 ;
        RECT 68.410 109.335 68.670 109.595 ;
        RECT 68.410 108.985 68.670 109.245 ;
        RECT 71.170 109.335 71.430 109.595 ;
        RECT 71.170 108.985 71.430 109.245 ;
        RECT 73.930 109.335 74.190 109.595 ;
        RECT 73.930 108.985 74.190 109.245 ;
        RECT 76.690 109.335 76.950 109.595 ;
        RECT 76.690 108.985 76.950 109.245 ;
        RECT 79.450 109.335 79.710 109.595 ;
        RECT 79.450 108.985 79.710 109.245 ;
        RECT 82.210 109.335 82.470 109.595 ;
        RECT 82.210 108.985 82.470 109.245 ;
        RECT 85.555 106.310 85.815 106.570 ;
        RECT 86.015 106.310 86.275 106.570 ;
        RECT 86.475 106.310 86.735 106.570 ;
        RECT 86.935 106.310 87.195 106.570 ;
        RECT 87.395 106.310 87.655 106.570 ;
        RECT 87.855 106.310 88.115 106.570 ;
        RECT 88.315 106.310 88.575 106.570 ;
        RECT 88.775 106.310 89.035 106.570 ;
        RECT 89.235 106.310 89.495 106.570 ;
        RECT 89.695 106.310 89.955 106.570 ;
        RECT 90.155 106.310 90.415 106.570 ;
        RECT 90.615 106.310 90.875 106.570 ;
        RECT 91.075 106.310 91.335 106.570 ;
        RECT 91.535 106.310 91.795 106.570 ;
        RECT 91.995 106.310 92.255 106.570 ;
        RECT 92.455 106.310 92.715 106.570 ;
        RECT 92.915 106.310 93.175 106.570 ;
        RECT 93.375 106.310 93.635 106.570 ;
        RECT 93.835 106.310 94.095 106.570 ;
        RECT 94.295 106.310 94.555 106.570 ;
        RECT 94.755 106.310 95.015 106.570 ;
        RECT 95.215 106.310 95.475 106.570 ;
        RECT 95.675 106.310 95.935 106.570 ;
        RECT 96.135 106.310 96.395 106.570 ;
        RECT 96.595 106.310 96.855 106.570 ;
        RECT 97.055 106.310 97.315 106.570 ;
        RECT 97.515 106.310 97.775 106.570 ;
        RECT 97.975 106.310 98.235 106.570 ;
        RECT 98.435 106.310 98.695 106.570 ;
        RECT 98.895 106.310 99.155 106.570 ;
        RECT 99.355 106.310 99.615 106.570 ;
        RECT 99.815 106.310 100.075 106.570 ;
        RECT 100.275 106.310 100.535 106.570 ;
        RECT 100.735 106.310 100.995 106.570 ;
        RECT 101.195 106.310 101.455 106.570 ;
        RECT 101.655 106.310 101.915 106.570 ;
        RECT 102.115 106.310 102.375 106.570 ;
        RECT 11.660 102.050 11.920 102.310 ;
        RECT 12.020 102.050 12.280 102.310 ;
        RECT 129.775 102.035 130.035 102.295 ;
        RECT 130.135 102.035 130.395 102.295 ;
        RECT 130.495 102.035 130.755 102.295 ;
        RECT 130.855 102.035 131.115 102.295 ;
        RECT 131.215 102.035 131.475 102.295 ;
        RECT 131.575 102.035 131.835 102.295 ;
        RECT 56.890 100.150 57.150 100.410 ;
        RECT 57.250 100.150 57.510 100.410 ;
        RECT 111.545 88.910 111.805 89.170 ;
        RECT 111.545 88.550 111.805 88.810 ;
        RECT 6.040 48.385 6.300 48.645 ;
        RECT 6.040 48.025 6.300 48.285 ;
        RECT 105.565 16.395 105.825 16.655 ;
        RECT 105.925 16.395 106.185 16.655 ;
        RECT 65.350 6.800 65.610 7.060 ;
        RECT 65.710 6.800 65.970 7.060 ;
        RECT 12.090 6.130 12.350 6.390 ;
        RECT 12.090 5.770 12.350 6.030 ;
      LAYER met2 ;
        RECT 21.430 108.930 21.810 110.420 ;
        RECT 24.190 108.930 24.570 110.420 ;
        RECT 26.950 108.930 27.330 110.420 ;
        RECT 29.710 108.930 30.090 110.420 ;
        RECT 32.470 108.930 32.850 110.420 ;
        RECT 35.230 108.930 35.610 110.420 ;
        RECT 37.990 108.930 38.370 110.420 ;
        RECT 40.750 108.930 41.130 110.420 ;
        RECT 43.510 108.930 43.890 110.420 ;
        RECT 46.270 108.930 46.650 110.420 ;
        RECT 49.030 108.930 49.410 110.420 ;
        RECT 51.790 108.930 52.170 110.420 ;
        RECT 54.550 108.930 54.930 110.420 ;
        RECT 57.310 108.930 57.690 110.420 ;
        RECT 60.070 108.930 60.450 110.420 ;
        RECT 62.830 108.930 63.210 110.420 ;
        RECT 65.590 108.930 65.970 110.420 ;
        RECT 68.350 108.930 68.730 110.420 ;
        RECT 71.110 108.930 71.490 110.420 ;
        RECT 73.870 108.930 74.250 110.420 ;
        RECT 76.630 108.930 77.010 110.420 ;
        RECT 79.390 108.930 79.770 110.420 ;
        RECT 82.150 108.930 82.530 110.420 ;
        RECT 84.955 105.700 102.975 107.180 ;
        RECT 11.130 101.520 12.810 102.840 ;
        RECT 13.235 102.345 17.915 103.025 ;
        RECT 129.245 101.505 132.365 102.825 ;
        RECT 56.360 99.620 58.040 100.940 ;
        RECT 58.500 100.495 63.180 101.175 ;
        RECT 111.015 88.020 112.335 89.700 ;
        RECT 111.835 82.880 112.515 87.560 ;
        RECT 5.295 49.610 5.975 54.290 ;
        RECT 5.510 47.495 6.830 49.175 ;
        RECT 99.920 15.665 104.600 16.345 ;
        RECT 105.035 15.865 106.715 17.185 ;
        RECT 11.270 7.410 11.950 12.090 ;
        RECT 11.560 5.240 12.880 6.920 ;
        RECT 59.710 6.095 64.390 6.775 ;
        RECT 64.820 6.270 66.500 7.590 ;
      LAYER via2 ;
        RECT 21.480 110.100 21.760 110.380 ;
        RECT 21.480 109.700 21.760 109.980 ;
        RECT 24.240 110.100 24.520 110.380 ;
        RECT 24.240 109.700 24.520 109.980 ;
        RECT 27.000 110.100 27.280 110.380 ;
        RECT 27.000 109.700 27.280 109.980 ;
        RECT 29.760 110.100 30.040 110.380 ;
        RECT 29.760 109.700 30.040 109.980 ;
        RECT 32.520 110.100 32.800 110.380 ;
        RECT 32.520 109.700 32.800 109.980 ;
        RECT 35.280 110.100 35.560 110.380 ;
        RECT 35.280 109.700 35.560 109.980 ;
        RECT 38.040 110.100 38.320 110.380 ;
        RECT 38.040 109.700 38.320 109.980 ;
        RECT 40.800 110.100 41.080 110.380 ;
        RECT 40.800 109.700 41.080 109.980 ;
        RECT 43.560 110.100 43.840 110.380 ;
        RECT 43.560 109.700 43.840 109.980 ;
        RECT 46.320 110.100 46.600 110.380 ;
        RECT 46.320 109.700 46.600 109.980 ;
        RECT 49.080 110.100 49.360 110.380 ;
        RECT 49.080 109.700 49.360 109.980 ;
        RECT 51.840 110.100 52.120 110.380 ;
        RECT 51.840 109.700 52.120 109.980 ;
        RECT 54.600 110.100 54.880 110.380 ;
        RECT 54.600 109.700 54.880 109.980 ;
        RECT 57.360 110.100 57.640 110.380 ;
        RECT 57.360 109.700 57.640 109.980 ;
        RECT 60.120 110.100 60.400 110.380 ;
        RECT 60.120 109.700 60.400 109.980 ;
        RECT 62.880 110.100 63.160 110.380 ;
        RECT 62.880 109.700 63.160 109.980 ;
        RECT 65.640 110.100 65.920 110.380 ;
        RECT 65.640 109.700 65.920 109.980 ;
        RECT 68.400 110.100 68.680 110.380 ;
        RECT 68.400 109.700 68.680 109.980 ;
        RECT 71.160 110.100 71.440 110.380 ;
        RECT 71.160 109.700 71.440 109.980 ;
        RECT 73.920 110.100 74.200 110.380 ;
        RECT 73.920 109.700 74.200 109.980 ;
        RECT 76.680 110.100 76.960 110.380 ;
        RECT 76.680 109.700 76.960 109.980 ;
        RECT 79.440 110.100 79.720 110.380 ;
        RECT 79.440 109.700 79.720 109.980 ;
        RECT 82.200 110.100 82.480 110.380 ;
        RECT 82.200 109.700 82.480 109.980 ;
        RECT 85.630 106.300 85.910 106.580 ;
        RECT 86.030 106.300 86.310 106.580 ;
        RECT 86.430 106.300 86.710 106.580 ;
        RECT 86.830 106.300 87.110 106.580 ;
        RECT 87.230 106.300 87.510 106.580 ;
        RECT 87.630 106.300 87.910 106.580 ;
        RECT 88.030 106.300 88.310 106.580 ;
        RECT 88.430 106.300 88.710 106.580 ;
        RECT 88.830 106.300 89.110 106.580 ;
        RECT 89.230 106.300 89.510 106.580 ;
        RECT 89.630 106.300 89.910 106.580 ;
        RECT 90.030 106.300 90.310 106.580 ;
        RECT 90.430 106.300 90.710 106.580 ;
        RECT 90.830 106.300 91.110 106.580 ;
        RECT 91.230 106.300 91.510 106.580 ;
        RECT 91.630 106.300 91.910 106.580 ;
        RECT 92.030 106.300 92.310 106.580 ;
        RECT 92.430 106.300 92.710 106.580 ;
        RECT 92.830 106.300 93.110 106.580 ;
        RECT 93.230 106.300 93.510 106.580 ;
        RECT 93.630 106.300 93.910 106.580 ;
        RECT 94.030 106.300 94.310 106.580 ;
        RECT 94.430 106.300 94.710 106.580 ;
        RECT 94.830 106.300 95.110 106.580 ;
        RECT 95.230 106.300 95.510 106.580 ;
        RECT 95.630 106.300 95.910 106.580 ;
        RECT 96.030 106.300 96.310 106.580 ;
        RECT 96.430 106.300 96.710 106.580 ;
        RECT 96.830 106.300 97.110 106.580 ;
        RECT 97.230 106.300 97.510 106.580 ;
        RECT 97.630 106.300 97.910 106.580 ;
        RECT 98.030 106.300 98.310 106.580 ;
        RECT 98.430 106.300 98.710 106.580 ;
        RECT 98.830 106.300 99.110 106.580 ;
        RECT 99.230 106.300 99.510 106.580 ;
        RECT 99.630 106.300 99.910 106.580 ;
        RECT 100.030 106.300 100.310 106.580 ;
        RECT 100.430 106.300 100.710 106.580 ;
        RECT 100.830 106.300 101.110 106.580 ;
        RECT 101.230 106.300 101.510 106.580 ;
        RECT 101.630 106.300 101.910 106.580 ;
        RECT 102.030 106.300 102.310 106.580 ;
        RECT 11.630 102.040 11.910 102.320 ;
        RECT 12.030 102.040 12.310 102.320 ;
        RECT 129.765 102.025 130.045 102.305 ;
        RECT 130.215 102.025 130.495 102.305 ;
        RECT 130.665 102.025 130.945 102.305 ;
        RECT 131.115 102.025 131.395 102.305 ;
        RECT 131.565 102.025 131.845 102.305 ;
        RECT 56.940 100.140 57.220 100.420 ;
        RECT 57.340 100.140 57.620 100.420 ;
        RECT 111.535 88.920 111.815 89.200 ;
        RECT 111.535 88.520 111.815 88.800 ;
        RECT 6.030 48.395 6.310 48.675 ;
        RECT 6.030 47.995 6.310 48.275 ;
        RECT 105.535 16.385 105.815 16.665 ;
        RECT 105.935 16.385 106.215 16.665 ;
        RECT 65.320 6.790 65.600 7.070 ;
        RECT 65.720 6.790 66.000 7.070 ;
        RECT 12.080 6.140 12.360 6.420 ;
        RECT 12.080 5.740 12.360 6.020 ;
      LAYER met3 ;
        RECT 10.690 109.040 82.530 110.425 ;
        RECT 138.730 109.040 157.320 111.520 ;
        RECT 10.690 105.580 157.320 109.040 ;
        RECT 10.690 99.620 83.670 105.580 ;
        RECT 111.355 90.140 157.320 105.580 ;
        RECT 3.000 46.230 14.740 54.365 ;
        RECT 3.000 4.200 20.790 46.230 ;
        RECT 109.910 25.070 157.320 90.140 ;
        RECT 99.815 7.585 157.320 25.070 ;
        RECT 59.425 4.200 157.320 7.585 ;
        RECT 3.000 0.000 157.320 4.200 ;
      LAYER via3 ;
        RECT 21.460 110.080 21.780 110.400 ;
        RECT 24.220 110.080 24.540 110.400 ;
        RECT 26.980 110.080 27.300 110.400 ;
        RECT 29.740 110.080 30.060 110.400 ;
        RECT 32.500 110.080 32.820 110.400 ;
        RECT 35.260 110.080 35.580 110.400 ;
        RECT 38.020 110.080 38.340 110.400 ;
        RECT 40.780 110.080 41.100 110.400 ;
        RECT 43.540 110.080 43.860 110.400 ;
        RECT 46.300 110.080 46.620 110.400 ;
        RECT 49.060 110.080 49.380 110.400 ;
        RECT 51.820 110.080 52.140 110.400 ;
        RECT 54.580 110.080 54.900 110.400 ;
        RECT 57.340 110.080 57.660 110.400 ;
        RECT 60.100 110.080 60.420 110.400 ;
        RECT 62.860 110.080 63.180 110.400 ;
        RECT 65.620 110.080 65.940 110.400 ;
        RECT 68.380 110.080 68.700 110.400 ;
        RECT 71.140 110.080 71.460 110.400 ;
        RECT 73.900 110.080 74.220 110.400 ;
        RECT 76.660 110.080 76.980 110.400 ;
        RECT 79.420 110.080 79.740 110.400 ;
        RECT 82.180 110.080 82.500 110.400 ;
        RECT 21.460 109.680 21.780 110.000 ;
        RECT 24.220 109.680 24.540 110.000 ;
        RECT 26.980 109.680 27.300 110.000 ;
        RECT 29.740 109.680 30.060 110.000 ;
        RECT 32.500 109.680 32.820 110.000 ;
        RECT 35.260 109.680 35.580 110.000 ;
        RECT 38.020 109.680 38.340 110.000 ;
        RECT 40.780 109.680 41.100 110.000 ;
        RECT 43.540 109.680 43.860 110.000 ;
        RECT 46.300 109.680 46.620 110.000 ;
        RECT 49.060 109.680 49.380 110.000 ;
        RECT 51.820 109.680 52.140 110.000 ;
        RECT 54.580 109.680 54.900 110.000 ;
        RECT 57.340 109.680 57.660 110.000 ;
        RECT 60.100 109.680 60.420 110.000 ;
        RECT 62.860 109.680 63.180 110.000 ;
        RECT 65.620 109.680 65.940 110.000 ;
        RECT 68.380 109.680 68.700 110.000 ;
        RECT 71.140 109.680 71.460 110.000 ;
        RECT 73.900 109.680 74.220 110.000 ;
        RECT 76.660 109.680 76.980 110.000 ;
        RECT 79.420 109.680 79.740 110.000 ;
        RECT 82.180 109.680 82.500 110.000 ;
        RECT 155.560 0.200 157.080 111.320 ;
      LAYER met4 ;
        RECT 21.470 110.425 21.770 111.520 ;
        RECT 24.230 110.425 24.530 111.520 ;
        RECT 26.990 110.425 27.290 111.520 ;
        RECT 29.750 110.425 30.050 111.520 ;
        RECT 32.510 110.425 32.810 111.520 ;
        RECT 35.270 110.425 35.570 111.520 ;
        RECT 38.030 110.425 38.330 111.520 ;
        RECT 40.790 110.425 41.090 111.520 ;
        RECT 43.550 110.425 43.850 111.520 ;
        RECT 46.310 110.425 46.610 111.520 ;
        RECT 49.070 110.425 49.370 111.520 ;
        RECT 51.830 110.425 52.130 111.520 ;
        RECT 54.590 110.425 54.890 111.520 ;
        RECT 57.350 110.425 57.650 111.520 ;
        RECT 60.110 110.425 60.410 111.520 ;
        RECT 62.870 110.425 63.170 111.520 ;
        RECT 65.630 110.425 65.930 111.520 ;
        RECT 68.390 110.425 68.690 111.520 ;
        RECT 71.150 110.425 71.450 111.520 ;
        RECT 73.910 110.425 74.210 111.520 ;
        RECT 76.670 110.425 76.970 111.520 ;
        RECT 79.430 110.425 79.730 111.520 ;
        RECT 82.190 110.425 82.490 111.520 ;
        RECT 21.430 109.650 21.810 110.425 ;
        RECT 24.190 109.650 24.570 110.425 ;
        RECT 26.950 109.650 27.330 110.425 ;
        RECT 29.710 109.650 30.090 110.425 ;
        RECT 32.470 109.650 32.850 110.425 ;
        RECT 35.230 109.650 35.610 110.425 ;
        RECT 37.990 109.650 38.370 110.425 ;
        RECT 40.750 109.650 41.130 110.425 ;
        RECT 43.510 109.650 43.890 110.425 ;
        RECT 46.270 109.650 46.650 110.425 ;
        RECT 49.030 109.650 49.410 110.425 ;
        RECT 51.790 109.650 52.170 110.425 ;
        RECT 54.550 109.650 54.930 110.425 ;
        RECT 57.310 109.650 57.690 110.425 ;
        RECT 60.070 109.650 60.450 110.425 ;
        RECT 62.830 109.650 63.210 110.425 ;
        RECT 65.590 109.650 65.970 110.425 ;
        RECT 68.350 109.650 68.730 110.425 ;
        RECT 71.110 109.650 71.490 110.425 ;
        RECT 73.870 109.650 74.250 110.425 ;
        RECT 76.630 109.650 77.010 110.425 ;
        RECT 79.390 109.650 79.770 110.425 ;
        RECT 82.150 109.650 82.530 110.425 ;
        RECT 155.320 0.000 157.320 111.520 ;
    END
  END VGND
  PIN clk
    PORT
      LAYER met1 ;
        RECT 134.595 108.930 134.965 109.650 ;
      LAYER via ;
        RECT 134.650 109.335 134.910 109.595 ;
        RECT 134.650 108.985 134.910 109.245 ;
      LAYER met2 ;
        RECT 134.590 108.930 134.970 110.420 ;
      LAYER via2 ;
        RECT 134.640 110.100 134.920 110.380 ;
        RECT 134.640 109.700 134.920 109.980 ;
      LAYER met3 ;
        RECT 134.590 109.650 134.970 110.425 ;
      LAYER via3 ;
        RECT 134.620 110.080 134.940 110.400 ;
        RECT 134.620 109.680 134.940 110.000 ;
      LAYER met4 ;
        RECT 134.630 110.425 134.930 111.520 ;
        RECT 134.590 109.650 134.970 110.425 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met1 ;
        RECT 137.355 108.930 137.725 109.650 ;
      LAYER via ;
        RECT 137.410 109.335 137.670 109.595 ;
        RECT 137.410 108.985 137.670 109.245 ;
      LAYER met2 ;
        RECT 137.350 108.930 137.730 110.420 ;
      LAYER via2 ;
        RECT 137.400 110.100 137.680 110.380 ;
        RECT 137.400 109.700 137.680 109.980 ;
      LAYER met3 ;
        RECT 137.350 109.650 137.730 110.425 ;
      LAYER via3 ;
        RECT 137.380 110.080 137.700 110.400 ;
        RECT 137.380 109.680 137.700 110.000 ;
      LAYER met4 ;
        RECT 137.390 110.425 137.690 111.520 ;
        RECT 137.350 109.650 137.730 110.425 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met1 ;
        RECT 131.835 108.930 132.205 109.650 ;
      LAYER via ;
        RECT 131.890 109.335 132.150 109.595 ;
        RECT 131.890 108.985 132.150 109.245 ;
      LAYER met2 ;
        RECT 131.830 108.930 132.210 110.420 ;
      LAYER via2 ;
        RECT 131.880 110.100 132.160 110.380 ;
        RECT 131.880 109.700 132.160 109.980 ;
      LAYER met3 ;
        RECT 131.830 109.650 132.210 110.425 ;
      LAYER via3 ;
        RECT 131.860 110.080 132.180 110.400 ;
        RECT 131.860 109.680 132.180 110.000 ;
      LAYER met4 ;
        RECT 131.870 110.425 132.170 111.520 ;
        RECT 131.830 109.650 132.210 110.425 ;
    END
  END rst_n
  PIN ui_in[0]
    PORT
      LAYER li1 ;
        RECT 129.710 103.260 131.890 103.610 ;
      LAYER mcon ;
        RECT 129.820 103.350 129.990 103.520 ;
        RECT 130.180 103.350 130.350 103.520 ;
        RECT 130.540 103.350 130.710 103.520 ;
        RECT 130.900 103.350 131.070 103.520 ;
        RECT 131.260 103.350 131.430 103.520 ;
        RECT 131.620 103.350 131.790 103.520 ;
      LAYER met1 ;
        RECT 129.075 108.930 129.445 109.650 ;
        RECT 129.075 108.630 130.060 108.930 ;
        RECT 129.760 103.860 130.060 108.630 ;
        RECT 129.755 103.310 131.860 103.860 ;
      LAYER via ;
        RECT 129.130 109.335 129.390 109.595 ;
        RECT 129.130 108.985 129.390 109.245 ;
      LAYER met2 ;
        RECT 129.070 108.930 129.450 110.420 ;
      LAYER via2 ;
        RECT 129.120 110.100 129.400 110.380 ;
        RECT 129.120 109.700 129.400 109.980 ;
      LAYER met3 ;
        RECT 129.070 109.650 129.450 110.425 ;
      LAYER via3 ;
        RECT 129.100 110.080 129.420 110.400 ;
        RECT 129.100 109.680 129.420 110.000 ;
      LAYER met4 ;
        RECT 129.110 110.425 129.410 111.520 ;
        RECT 129.070 109.650 129.450 110.425 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER li1 ;
        RECT 127.225 104.530 129.405 104.880 ;
      LAYER mcon ;
        RECT 127.335 104.620 127.505 104.790 ;
        RECT 127.695 104.620 127.865 104.790 ;
        RECT 128.055 104.620 128.225 104.790 ;
        RECT 128.415 104.620 128.585 104.790 ;
        RECT 128.775 104.620 128.945 104.790 ;
        RECT 129.135 104.620 129.305 104.790 ;
      LAYER met1 ;
        RECT 126.315 108.930 126.685 109.650 ;
        RECT 126.315 108.630 127.570 108.930 ;
        RECT 127.275 105.130 127.575 108.630 ;
        RECT 127.270 104.580 129.375 105.130 ;
      LAYER via ;
        RECT 126.370 109.335 126.630 109.595 ;
        RECT 126.370 108.985 126.630 109.245 ;
      LAYER met2 ;
        RECT 126.310 108.930 126.690 110.420 ;
      LAYER via2 ;
        RECT 126.360 110.100 126.640 110.380 ;
        RECT 126.360 109.700 126.640 109.980 ;
      LAYER met3 ;
        RECT 126.310 109.650 126.690 110.425 ;
      LAYER via3 ;
        RECT 126.340 110.080 126.660 110.400 ;
        RECT 126.340 109.680 126.660 110.000 ;
      LAYER met4 ;
        RECT 126.350 110.425 126.650 111.520 ;
        RECT 126.310 109.650 126.690 110.425 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER li1 ;
        RECT 124.740 105.800 126.920 106.150 ;
      LAYER mcon ;
        RECT 124.850 105.890 125.020 106.060 ;
        RECT 125.210 105.890 125.380 106.060 ;
        RECT 125.570 105.890 125.740 106.060 ;
        RECT 125.930 105.890 126.100 106.060 ;
        RECT 126.290 105.890 126.460 106.060 ;
        RECT 126.650 105.890 126.820 106.060 ;
      LAYER met1 ;
        RECT 123.555 108.930 123.925 109.650 ;
        RECT 123.555 108.630 125.090 108.930 ;
        RECT 124.790 106.400 125.090 108.630 ;
        RECT 124.785 105.850 126.890 106.400 ;
      LAYER via ;
        RECT 123.610 109.335 123.870 109.595 ;
        RECT 123.610 108.985 123.870 109.245 ;
      LAYER met2 ;
        RECT 123.550 108.930 123.930 110.420 ;
      LAYER via2 ;
        RECT 123.600 110.100 123.880 110.380 ;
        RECT 123.600 109.700 123.880 109.980 ;
      LAYER met3 ;
        RECT 123.550 109.650 123.930 110.425 ;
      LAYER via3 ;
        RECT 123.580 110.080 123.900 110.400 ;
        RECT 123.580 109.680 123.900 110.000 ;
      LAYER met4 ;
        RECT 123.590 110.425 123.890 111.520 ;
        RECT 123.550 109.650 123.930 110.425 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER li1 ;
        RECT 122.255 107.070 124.435 107.420 ;
      LAYER mcon ;
        RECT 122.365 107.160 122.535 107.330 ;
        RECT 122.725 107.160 122.895 107.330 ;
        RECT 123.085 107.160 123.255 107.330 ;
        RECT 123.445 107.160 123.615 107.330 ;
        RECT 123.805 107.160 123.975 107.330 ;
        RECT 124.165 107.160 124.335 107.330 ;
      LAYER met1 ;
        RECT 120.795 108.930 121.165 109.650 ;
        RECT 120.795 108.630 122.605 108.930 ;
        RECT 122.305 107.670 122.605 108.630 ;
        RECT 122.300 107.120 124.405 107.670 ;
      LAYER via ;
        RECT 120.850 109.335 121.110 109.595 ;
        RECT 120.850 108.985 121.110 109.245 ;
      LAYER met2 ;
        RECT 120.790 108.930 121.170 110.420 ;
      LAYER via2 ;
        RECT 120.840 110.100 121.120 110.380 ;
        RECT 120.840 109.700 121.120 109.980 ;
      LAYER met3 ;
        RECT 120.790 109.650 121.170 110.425 ;
      LAYER via3 ;
        RECT 120.820 110.080 121.140 110.400 ;
        RECT 120.820 109.680 121.140 110.000 ;
      LAYER met4 ;
        RECT 120.830 110.425 121.130 111.520 ;
        RECT 120.790 109.650 121.170 110.425 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER li1 ;
        RECT 114.395 107.070 116.575 107.420 ;
      LAYER mcon ;
        RECT 114.490 107.160 114.660 107.330 ;
        RECT 114.850 107.160 115.020 107.330 ;
        RECT 115.210 107.160 115.380 107.330 ;
        RECT 115.570 107.160 115.740 107.330 ;
        RECT 115.930 107.160 116.100 107.330 ;
        RECT 116.290 107.160 116.460 107.330 ;
      LAYER met1 ;
        RECT 118.035 108.930 118.405 109.650 ;
        RECT 116.230 108.630 118.405 108.930 ;
        RECT 116.230 107.670 116.530 108.630 ;
        RECT 114.425 107.120 116.530 107.670 ;
      LAYER via ;
        RECT 118.090 109.335 118.350 109.595 ;
        RECT 118.090 108.985 118.350 109.245 ;
      LAYER met2 ;
        RECT 118.030 108.930 118.410 110.420 ;
      LAYER via2 ;
        RECT 118.080 110.100 118.360 110.380 ;
        RECT 118.080 109.700 118.360 109.980 ;
      LAYER met3 ;
        RECT 118.030 109.650 118.410 110.425 ;
      LAYER via3 ;
        RECT 118.060 110.080 118.380 110.400 ;
        RECT 118.060 109.680 118.380 110.000 ;
      LAYER met4 ;
        RECT 118.070 110.425 118.370 111.520 ;
        RECT 118.030 109.650 118.410 110.425 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER li1 ;
        RECT 111.910 105.800 114.090 106.150 ;
      LAYER mcon ;
        RECT 112.005 105.890 112.175 106.060 ;
        RECT 112.365 105.890 112.535 106.060 ;
        RECT 112.725 105.890 112.895 106.060 ;
        RECT 113.085 105.890 113.255 106.060 ;
        RECT 113.445 105.890 113.615 106.060 ;
        RECT 113.805 105.890 113.975 106.060 ;
      LAYER met1 ;
        RECT 115.275 108.930 115.645 109.650 ;
        RECT 113.745 108.630 115.645 108.930 ;
        RECT 113.745 106.400 114.045 108.630 ;
        RECT 111.940 105.850 114.045 106.400 ;
      LAYER via ;
        RECT 115.330 109.335 115.590 109.595 ;
        RECT 115.330 108.985 115.590 109.245 ;
      LAYER met2 ;
        RECT 115.270 108.930 115.650 110.420 ;
      LAYER via2 ;
        RECT 115.320 110.100 115.600 110.380 ;
        RECT 115.320 109.700 115.600 109.980 ;
      LAYER met3 ;
        RECT 115.270 109.650 115.650 110.425 ;
      LAYER via3 ;
        RECT 115.300 110.080 115.620 110.400 ;
        RECT 115.300 109.680 115.620 110.000 ;
      LAYER met4 ;
        RECT 115.310 110.425 115.610 111.520 ;
        RECT 115.270 109.650 115.650 110.425 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER li1 ;
        RECT 109.425 104.530 111.605 104.880 ;
      LAYER mcon ;
        RECT 109.520 104.620 109.690 104.790 ;
        RECT 109.880 104.620 110.050 104.790 ;
        RECT 110.240 104.620 110.410 104.790 ;
        RECT 110.600 104.620 110.770 104.790 ;
        RECT 110.960 104.620 111.130 104.790 ;
        RECT 111.320 104.620 111.490 104.790 ;
      LAYER met1 ;
        RECT 112.515 108.930 112.885 109.650 ;
        RECT 111.260 108.630 112.885 108.930 ;
        RECT 111.260 105.130 111.560 108.630 ;
        RECT 109.455 104.580 111.560 105.130 ;
      LAYER via ;
        RECT 112.570 109.335 112.830 109.595 ;
        RECT 112.570 108.985 112.830 109.245 ;
      LAYER met2 ;
        RECT 112.510 108.930 112.890 110.420 ;
      LAYER via2 ;
        RECT 112.560 110.100 112.840 110.380 ;
        RECT 112.560 109.700 112.840 109.980 ;
      LAYER met3 ;
        RECT 112.510 109.650 112.890 110.425 ;
      LAYER via3 ;
        RECT 112.540 110.080 112.860 110.400 ;
        RECT 112.540 109.680 112.860 110.000 ;
      LAYER met4 ;
        RECT 112.550 110.425 112.850 111.520 ;
        RECT 112.510 109.650 112.890 110.425 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER li1 ;
        RECT 106.940 103.260 109.120 103.610 ;
      LAYER mcon ;
        RECT 107.035 103.350 107.205 103.520 ;
        RECT 107.395 103.350 107.565 103.520 ;
        RECT 107.755 103.350 107.925 103.520 ;
        RECT 108.115 103.350 108.285 103.520 ;
        RECT 108.475 103.350 108.645 103.520 ;
        RECT 108.835 103.350 109.005 103.520 ;
      LAYER met1 ;
        RECT 109.755 108.930 110.125 109.650 ;
        RECT 108.775 108.630 110.125 108.930 ;
        RECT 108.775 103.860 109.075 108.630 ;
        RECT 106.970 103.310 109.075 103.860 ;
      LAYER via ;
        RECT 109.810 109.335 110.070 109.595 ;
        RECT 109.810 108.985 110.070 109.245 ;
      LAYER met2 ;
        RECT 109.750 108.930 110.130 110.420 ;
      LAYER via2 ;
        RECT 109.800 110.100 110.080 110.380 ;
        RECT 109.800 109.700 110.080 109.980 ;
      LAYER met3 ;
        RECT 109.750 109.650 110.130 110.425 ;
      LAYER via3 ;
        RECT 109.780 110.080 110.100 110.400 ;
        RECT 109.780 109.680 110.100 110.000 ;
      LAYER met4 ;
        RECT 109.790 110.425 110.090 111.520 ;
        RECT 109.750 109.650 110.130 110.425 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met1 ;
        RECT 106.995 108.930 107.365 109.650 ;
      LAYER via ;
        RECT 107.050 109.335 107.310 109.595 ;
        RECT 107.050 108.985 107.310 109.245 ;
      LAYER met2 ;
        RECT 106.990 108.930 107.370 110.420 ;
      LAYER via2 ;
        RECT 107.040 110.100 107.320 110.380 ;
        RECT 107.040 109.700 107.320 109.980 ;
      LAYER met3 ;
        RECT 106.990 109.650 107.370 110.425 ;
      LAYER via3 ;
        RECT 107.020 110.080 107.340 110.400 ;
        RECT 107.020 109.680 107.340 110.000 ;
      LAYER met4 ;
        RECT 107.030 110.425 107.330 111.520 ;
        RECT 106.990 109.650 107.370 110.425 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met1 ;
        RECT 104.235 108.930 104.605 109.650 ;
      LAYER via ;
        RECT 104.290 109.335 104.550 109.595 ;
        RECT 104.290 108.985 104.550 109.245 ;
      LAYER met2 ;
        RECT 104.230 108.930 104.610 110.420 ;
      LAYER via2 ;
        RECT 104.280 110.100 104.560 110.380 ;
        RECT 104.280 109.700 104.560 109.980 ;
      LAYER met3 ;
        RECT 104.230 109.650 104.610 110.425 ;
      LAYER via3 ;
        RECT 104.260 110.080 104.580 110.400 ;
        RECT 104.260 109.680 104.580 110.000 ;
      LAYER met4 ;
        RECT 104.270 110.425 104.570 111.520 ;
        RECT 104.230 109.650 104.610 110.425 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met1 ;
        RECT 101.475 108.930 101.845 109.650 ;
      LAYER via ;
        RECT 101.530 109.335 101.790 109.595 ;
        RECT 101.530 108.985 101.790 109.245 ;
      LAYER met2 ;
        RECT 101.470 108.930 101.850 110.420 ;
      LAYER via2 ;
        RECT 101.520 110.100 101.800 110.380 ;
        RECT 101.520 109.700 101.800 109.980 ;
      LAYER met3 ;
        RECT 101.470 109.650 101.850 110.425 ;
      LAYER via3 ;
        RECT 101.500 110.080 101.820 110.400 ;
        RECT 101.500 109.680 101.820 110.000 ;
      LAYER met4 ;
        RECT 101.510 110.425 101.810 111.520 ;
        RECT 101.470 109.650 101.850 110.425 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met1 ;
        RECT 98.715 108.930 99.085 109.650 ;
      LAYER via ;
        RECT 98.770 109.335 99.030 109.595 ;
        RECT 98.770 108.985 99.030 109.245 ;
      LAYER met2 ;
        RECT 98.710 108.930 99.090 110.420 ;
      LAYER via2 ;
        RECT 98.760 110.100 99.040 110.380 ;
        RECT 98.760 109.700 99.040 109.980 ;
      LAYER met3 ;
        RECT 98.710 109.650 99.090 110.425 ;
      LAYER via3 ;
        RECT 98.740 110.080 99.060 110.400 ;
        RECT 98.740 109.680 99.060 110.000 ;
      LAYER met4 ;
        RECT 98.750 110.425 99.050 111.520 ;
        RECT 98.710 109.650 99.090 110.425 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met1 ;
        RECT 95.955 108.930 96.325 109.650 ;
      LAYER via ;
        RECT 96.010 109.335 96.270 109.595 ;
        RECT 96.010 108.985 96.270 109.245 ;
      LAYER met2 ;
        RECT 95.950 108.930 96.330 110.420 ;
      LAYER via2 ;
        RECT 96.000 110.100 96.280 110.380 ;
        RECT 96.000 109.700 96.280 109.980 ;
      LAYER met3 ;
        RECT 95.950 109.650 96.330 110.425 ;
      LAYER via3 ;
        RECT 95.980 110.080 96.300 110.400 ;
        RECT 95.980 109.680 96.300 110.000 ;
      LAYER met4 ;
        RECT 95.990 110.425 96.290 111.520 ;
        RECT 95.950 109.650 96.330 110.425 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met1 ;
        RECT 93.195 108.930 93.565 109.650 ;
      LAYER via ;
        RECT 93.250 109.335 93.510 109.595 ;
        RECT 93.250 108.985 93.510 109.245 ;
      LAYER met2 ;
        RECT 93.190 108.930 93.570 110.420 ;
      LAYER via2 ;
        RECT 93.240 110.100 93.520 110.380 ;
        RECT 93.240 109.700 93.520 109.980 ;
      LAYER met3 ;
        RECT 93.190 109.650 93.570 110.425 ;
      LAYER via3 ;
        RECT 93.220 110.080 93.540 110.400 ;
        RECT 93.220 109.680 93.540 110.000 ;
      LAYER met4 ;
        RECT 93.230 110.425 93.530 111.520 ;
        RECT 93.190 109.650 93.570 110.425 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met1 ;
        RECT 90.435 108.930 90.805 109.650 ;
      LAYER via ;
        RECT 90.490 109.335 90.750 109.595 ;
        RECT 90.490 108.985 90.750 109.245 ;
      LAYER met2 ;
        RECT 90.430 108.930 90.810 110.420 ;
      LAYER via2 ;
        RECT 90.480 110.100 90.760 110.380 ;
        RECT 90.480 109.700 90.760 109.980 ;
      LAYER met3 ;
        RECT 90.430 109.650 90.810 110.425 ;
      LAYER via3 ;
        RECT 90.460 110.080 90.780 110.400 ;
        RECT 90.460 109.680 90.780 110.000 ;
      LAYER met4 ;
        RECT 90.470 110.425 90.770 111.520 ;
        RECT 90.430 109.650 90.810 110.425 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met1 ;
        RECT 87.675 108.930 88.045 109.650 ;
      LAYER via ;
        RECT 87.730 109.335 87.990 109.595 ;
        RECT 87.730 108.985 87.990 109.245 ;
      LAYER met2 ;
        RECT 87.670 108.930 88.050 110.420 ;
      LAYER via2 ;
        RECT 87.720 110.100 88.000 110.380 ;
        RECT 87.720 109.700 88.000 109.980 ;
      LAYER met3 ;
        RECT 87.670 109.650 88.050 110.425 ;
      LAYER via3 ;
        RECT 87.700 110.080 88.020 110.400 ;
        RECT 87.700 109.680 88.020 110.000 ;
      LAYER met4 ;
        RECT 87.710 110.425 88.010 111.520 ;
        RECT 87.670 109.650 88.050 110.425 ;
    END
  END uio_in[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER li1 ;
        RECT 90.610 106.180 90.780 106.185 ;
        RECT 91.450 106.180 91.620 106.185 ;
        RECT 92.290 106.180 92.540 106.185 ;
        RECT 85.540 105.705 85.815 106.075 ;
        RECT 86.330 105.705 86.660 106.180 ;
        RECT 87.170 105.705 87.500 106.180 ;
        RECT 88.010 105.705 88.340 106.180 ;
        RECT 88.850 105.705 89.180 106.180 ;
        RECT 89.690 105.705 90.020 106.180 ;
        RECT 90.530 105.705 90.860 106.180 ;
        RECT 91.370 105.705 91.700 106.180 ;
        RECT 92.210 105.705 92.540 106.180 ;
        RECT 85.540 105.535 92.540 105.705 ;
        RECT 85.540 104.995 85.920 105.535 ;
        RECT 85.540 104.825 92.540 104.995 ;
        RECT 85.540 104.080 85.815 104.825 ;
        RECT 86.330 103.975 86.660 104.825 ;
        RECT 87.170 103.975 87.500 104.825 ;
        RECT 88.010 103.975 88.340 104.825 ;
        RECT 88.850 103.975 89.180 104.825 ;
        RECT 89.690 103.975 90.020 104.825 ;
        RECT 90.530 103.975 90.860 104.825 ;
        RECT 91.370 103.975 91.700 104.825 ;
        RECT 92.210 103.975 92.540 104.825 ;
      LAYER mcon ;
        RECT 85.595 105.860 85.765 106.030 ;
        RECT 85.595 105.430 85.765 105.600 ;
        RECT 85.595 104.995 85.765 105.165 ;
        RECT 85.595 104.560 85.765 104.730 ;
        RECT 85.595 104.130 85.765 104.300 ;
      LAYER met1 ;
        RECT 84.915 106.060 85.285 109.650 ;
        RECT 84.915 104.100 85.815 106.060 ;
      LAYER via ;
        RECT 84.970 109.335 85.230 109.595 ;
        RECT 84.970 108.985 85.230 109.245 ;
      LAYER met2 ;
        RECT 84.910 108.930 85.290 110.420 ;
      LAYER via2 ;
        RECT 84.960 110.100 85.240 110.380 ;
        RECT 84.960 109.700 85.240 109.980 ;
      LAYER met3 ;
        RECT 84.910 109.650 85.290 110.425 ;
      LAYER via3 ;
        RECT 84.940 110.080 85.260 110.400 ;
        RECT 84.940 109.680 85.260 110.000 ;
      LAYER met4 ;
        RECT 84.950 110.425 85.250 111.520 ;
        RECT 84.910 109.650 85.290 110.425 ;
    END
  END uo_out[0]
  PIN VPWR
    ANTENNADIFFAREA 661.659058 ;
    PORT
      LAYER nwell ;
        RECT 10.830 98.335 11.420 98.340 ;
        RECT 41.680 98.335 51.930 98.340 ;
        RECT 10.830 90.365 51.930 98.335 ;
        RECT 56.060 96.435 56.650 96.440 ;
        RECT 86.910 96.435 97.160 96.440 ;
        RECT 56.060 88.465 97.160 96.435 ;
        RECT 99.860 89.410 107.835 90.000 ;
        RECT 10.010 78.045 17.985 88.295 ;
        RECT 10.015 47.785 17.985 78.045 ;
        RECT 99.860 59.150 107.830 89.410 ;
        RECT 99.860 48.900 107.835 59.150 ;
        RECT 10.010 47.195 17.985 47.785 ;
        RECT 16.060 35.790 24.035 46.040 ;
        RECT 16.065 5.530 24.035 35.790 ;
        RECT 65.915 20.370 107.015 28.340 ;
        RECT 65.915 20.365 76.165 20.370 ;
        RECT 106.425 20.365 107.015 20.370 ;
        RECT 25.700 10.775 66.800 18.745 ;
        RECT 25.700 10.770 35.950 10.775 ;
        RECT 66.210 10.770 66.800 10.775 ;
        RECT 16.060 4.940 24.035 5.530 ;
      LAYER li1 ;
        RECT 85.990 103.805 86.160 104.605 ;
        RECT 86.830 103.805 87.000 104.605 ;
        RECT 87.670 103.805 87.840 104.605 ;
        RECT 88.510 103.805 88.680 104.605 ;
        RECT 89.350 103.805 89.520 104.605 ;
        RECT 90.190 103.805 90.360 104.605 ;
        RECT 91.030 103.805 91.200 104.605 ;
        RECT 91.870 103.805 92.040 104.605 ;
        RECT 92.710 103.805 92.880 104.605 ;
        RECT 93.550 103.805 93.720 104.605 ;
        RECT 94.390 103.805 94.560 104.605 ;
        RECT 95.230 103.805 95.400 104.995 ;
        RECT 96.050 103.805 96.380 104.955 ;
        RECT 96.890 103.805 97.220 104.605 ;
        RECT 97.730 103.805 98.060 104.605 ;
        RECT 98.570 103.805 98.900 104.605 ;
        RECT 99.490 103.805 99.660 104.605 ;
        RECT 100.330 103.805 100.500 104.605 ;
        RECT 101.620 103.805 101.950 104.565 ;
        RECT 85.455 103.635 102.475 103.805 ;
        RECT 107.190 101.990 109.370 102.340 ;
        RECT 11.585 92.060 51.515 92.950 ;
        RECT 11.585 90.885 51.515 91.775 ;
        RECT 56.815 90.160 96.745 91.050 ;
        RECT 56.815 88.985 96.745 89.875 ;
        RECT 15.400 47.950 16.290 87.880 ;
        RECT 16.575 47.950 17.465 87.880 ;
        RECT 100.380 49.315 101.270 89.245 ;
        RECT 101.555 49.315 102.445 89.245 ;
        RECT 21.450 5.695 22.340 45.625 ;
        RECT 22.625 5.695 23.515 45.625 ;
        RECT 66.330 26.930 106.260 27.820 ;
        RECT 66.330 25.755 106.260 26.645 ;
        RECT 26.115 17.335 66.045 18.225 ;
        RECT 26.115 16.160 66.045 17.050 ;
      LAYER mcon ;
        RECT 85.600 103.635 85.770 103.805 ;
        RECT 86.060 103.635 86.230 103.805 ;
        RECT 86.520 103.635 86.690 103.805 ;
        RECT 86.980 103.635 87.150 103.805 ;
        RECT 87.440 103.635 87.610 103.805 ;
        RECT 87.900 103.635 88.070 103.805 ;
        RECT 88.360 103.635 88.530 103.805 ;
        RECT 88.820 103.635 88.990 103.805 ;
        RECT 89.280 103.635 89.450 103.805 ;
        RECT 89.740 103.635 89.910 103.805 ;
        RECT 90.200 103.635 90.370 103.805 ;
        RECT 90.660 103.635 90.830 103.805 ;
        RECT 91.120 103.635 91.290 103.805 ;
        RECT 91.580 103.635 91.750 103.805 ;
        RECT 92.040 103.635 92.210 103.805 ;
        RECT 92.500 103.635 92.670 103.805 ;
        RECT 92.960 103.635 93.130 103.805 ;
        RECT 93.420 103.635 93.590 103.805 ;
        RECT 93.880 103.635 94.050 103.805 ;
        RECT 94.340 103.635 94.510 103.805 ;
        RECT 94.800 103.635 94.970 103.805 ;
        RECT 95.260 103.635 95.430 103.805 ;
        RECT 95.720 103.635 95.890 103.805 ;
        RECT 96.180 103.635 96.350 103.805 ;
        RECT 96.640 103.635 96.810 103.805 ;
        RECT 97.100 103.635 97.270 103.805 ;
        RECT 97.560 103.635 97.730 103.805 ;
        RECT 98.020 103.635 98.190 103.805 ;
        RECT 98.480 103.635 98.650 103.805 ;
        RECT 98.940 103.635 99.110 103.805 ;
        RECT 99.400 103.635 99.570 103.805 ;
        RECT 99.860 103.635 100.030 103.805 ;
        RECT 100.320 103.635 100.490 103.805 ;
        RECT 100.780 103.635 100.950 103.805 ;
        RECT 101.240 103.635 101.410 103.805 ;
        RECT 101.700 103.635 101.870 103.805 ;
        RECT 102.160 103.635 102.330 103.805 ;
        RECT 107.285 102.080 107.455 102.250 ;
        RECT 107.645 102.080 107.815 102.250 ;
        RECT 108.005 102.080 108.175 102.250 ;
        RECT 108.365 102.080 108.535 102.250 ;
        RECT 108.725 102.080 108.895 102.250 ;
        RECT 109.085 102.080 109.255 102.250 ;
        RECT 11.665 92.060 51.435 92.950 ;
        RECT 11.665 90.885 51.435 91.775 ;
        RECT 56.895 90.160 96.665 91.050 ;
        RECT 56.895 88.985 96.665 89.875 ;
        RECT 15.400 48.030 16.290 87.800 ;
        RECT 16.575 48.030 17.465 87.800 ;
        RECT 100.380 49.395 101.270 89.165 ;
        RECT 101.555 49.395 102.445 89.165 ;
        RECT 21.450 5.775 22.340 45.545 ;
        RECT 22.625 5.775 23.515 45.545 ;
        RECT 66.410 26.930 106.180 27.820 ;
        RECT 66.410 25.755 106.180 26.645 ;
        RECT 26.195 17.335 65.965 18.225 ;
        RECT 26.195 16.160 65.965 17.050 ;
      LAYER met1 ;
        RECT 85.455 103.480 102.475 103.960 ;
        RECT 91.300 102.095 91.560 102.355 ;
        RECT 91.700 102.095 91.960 102.355 ;
        RECT 92.100 102.095 92.360 102.355 ;
        RECT 92.500 102.095 92.760 102.355 ;
        RECT 92.900 102.095 93.160 102.355 ;
        RECT 93.300 102.095 93.560 102.355 ;
        RECT 93.700 102.095 93.960 102.355 ;
        RECT 94.100 102.095 94.360 102.355 ;
        RECT 94.500 102.095 94.760 102.355 ;
        RECT 94.900 102.095 95.160 102.355 ;
        RECT 95.300 102.095 95.560 102.355 ;
        RECT 95.700 102.095 95.960 102.355 ;
        RECT 107.210 102.005 109.330 102.325 ;
        RECT 91.300 101.695 91.560 101.955 ;
        RECT 91.700 101.695 91.960 101.955 ;
        RECT 92.100 101.695 92.360 101.955 ;
        RECT 92.500 101.695 92.760 101.955 ;
        RECT 92.900 101.695 93.160 101.955 ;
        RECT 93.300 101.695 93.560 101.955 ;
        RECT 93.700 101.695 93.960 101.955 ;
        RECT 94.100 101.695 94.360 101.955 ;
        RECT 94.500 101.695 94.760 101.955 ;
        RECT 94.900 101.695 95.160 101.955 ;
        RECT 95.300 101.695 95.560 101.955 ;
        RECT 95.700 101.695 95.960 101.955 ;
        RECT 11.605 91.775 51.495 92.980 ;
        RECT 11.585 90.840 51.515 91.775 ;
        RECT 56.835 89.875 96.725 91.080 ;
        RECT 56.815 88.940 96.745 89.875 ;
        RECT 100.335 89.225 101.270 89.245 ;
        RECT 16.575 87.860 17.510 87.880 ;
        RECT 15.370 47.970 17.510 87.860 ;
        RECT 100.335 49.335 102.475 89.225 ;
        RECT 100.335 49.315 101.270 49.335 ;
        RECT 16.575 47.950 17.510 47.970 ;
        RECT 22.625 45.605 23.560 45.625 ;
        RECT 21.420 5.715 23.560 45.605 ;
        RECT 66.330 26.930 106.260 27.865 ;
        RECT 66.350 25.725 106.240 26.930 ;
        RECT 26.115 17.335 66.045 18.270 ;
        RECT 26.135 16.130 66.025 17.335 ;
        RECT 22.625 5.695 23.560 5.715 ;
      LAYER via ;
        RECT 85.555 103.590 85.815 103.850 ;
        RECT 86.015 103.590 86.275 103.850 ;
        RECT 86.475 103.590 86.735 103.850 ;
        RECT 86.935 103.590 87.195 103.850 ;
        RECT 87.395 103.590 87.655 103.850 ;
        RECT 87.855 103.590 88.115 103.850 ;
        RECT 88.315 103.590 88.575 103.850 ;
        RECT 88.775 103.590 89.035 103.850 ;
        RECT 89.235 103.590 89.495 103.850 ;
        RECT 89.695 103.590 89.955 103.850 ;
        RECT 90.155 103.590 90.415 103.850 ;
        RECT 90.615 103.590 90.875 103.850 ;
        RECT 91.075 103.590 91.335 103.850 ;
        RECT 91.535 103.590 91.795 103.850 ;
        RECT 91.995 103.590 92.255 103.850 ;
        RECT 92.455 103.590 92.715 103.850 ;
        RECT 92.915 103.590 93.175 103.850 ;
        RECT 93.375 103.590 93.635 103.850 ;
        RECT 93.835 103.590 94.095 103.850 ;
        RECT 94.295 103.590 94.555 103.850 ;
        RECT 94.755 103.590 95.015 103.850 ;
        RECT 95.215 103.590 95.475 103.850 ;
        RECT 95.675 103.590 95.935 103.850 ;
        RECT 96.135 103.590 96.395 103.850 ;
        RECT 96.595 103.590 96.855 103.850 ;
        RECT 97.055 103.590 97.315 103.850 ;
        RECT 97.515 103.590 97.775 103.850 ;
        RECT 97.975 103.590 98.235 103.850 ;
        RECT 98.435 103.590 98.695 103.850 ;
        RECT 98.895 103.590 99.155 103.850 ;
        RECT 99.355 103.590 99.615 103.850 ;
        RECT 99.815 103.590 100.075 103.850 ;
        RECT 100.275 103.590 100.535 103.850 ;
        RECT 100.735 103.590 100.995 103.850 ;
        RECT 101.195 103.590 101.455 103.850 ;
        RECT 101.655 103.590 101.915 103.850 ;
        RECT 102.115 103.590 102.375 103.850 ;
        RECT 107.240 102.035 107.500 102.295 ;
        RECT 107.600 102.035 107.860 102.295 ;
        RECT 107.960 102.035 108.220 102.295 ;
        RECT 108.320 102.035 108.580 102.295 ;
        RECT 108.680 102.035 108.940 102.295 ;
        RECT 109.040 102.035 109.300 102.295 ;
        RECT 11.620 91.560 11.880 91.820 ;
        RECT 11.980 91.560 12.240 91.820 ;
        RECT 12.340 91.560 12.600 91.820 ;
        RECT 12.700 91.560 12.960 91.820 ;
        RECT 13.060 91.560 13.320 91.820 ;
        RECT 13.420 91.560 13.680 91.820 ;
        RECT 13.780 91.560 14.040 91.820 ;
        RECT 14.140 91.560 14.400 91.820 ;
        RECT 14.500 91.560 14.760 91.820 ;
        RECT 14.860 91.560 15.120 91.820 ;
        RECT 15.220 91.560 15.480 91.820 ;
        RECT 15.580 91.560 15.840 91.820 ;
        RECT 15.940 91.560 16.200 91.820 ;
        RECT 16.300 91.560 16.560 91.820 ;
        RECT 16.660 91.560 16.920 91.820 ;
        RECT 17.020 91.560 17.280 91.820 ;
        RECT 17.380 91.560 17.640 91.820 ;
        RECT 17.740 91.560 18.000 91.820 ;
        RECT 18.100 91.560 18.360 91.820 ;
        RECT 18.460 91.560 18.720 91.820 ;
        RECT 18.820 91.560 19.080 91.820 ;
        RECT 19.180 91.560 19.440 91.820 ;
        RECT 19.540 91.560 19.800 91.820 ;
        RECT 19.900 91.560 20.160 91.820 ;
        RECT 20.260 91.560 20.520 91.820 ;
        RECT 20.620 91.560 20.880 91.820 ;
        RECT 20.980 91.560 21.240 91.820 ;
        RECT 21.340 91.560 21.600 91.820 ;
        RECT 21.700 91.560 21.960 91.820 ;
        RECT 22.060 91.560 22.320 91.820 ;
        RECT 22.420 91.560 22.680 91.820 ;
        RECT 22.780 91.560 23.040 91.820 ;
        RECT 23.140 91.560 23.400 91.820 ;
        RECT 23.500 91.560 23.760 91.820 ;
        RECT 23.860 91.560 24.120 91.820 ;
        RECT 24.220 91.560 24.480 91.820 ;
        RECT 24.580 91.560 24.840 91.820 ;
        RECT 24.940 91.560 25.200 91.820 ;
        RECT 25.300 91.560 25.560 91.820 ;
        RECT 25.660 91.560 25.920 91.820 ;
        RECT 26.020 91.560 26.280 91.820 ;
        RECT 26.380 91.560 26.640 91.820 ;
        RECT 26.740 91.560 27.000 91.820 ;
        RECT 27.100 91.560 27.360 91.820 ;
        RECT 27.460 91.560 27.720 91.820 ;
        RECT 27.820 91.560 28.080 91.820 ;
        RECT 28.180 91.560 28.440 91.820 ;
        RECT 28.540 91.560 28.800 91.820 ;
        RECT 28.900 91.560 29.160 91.820 ;
        RECT 29.260 91.560 29.520 91.820 ;
        RECT 29.620 91.560 29.880 91.820 ;
        RECT 29.980 91.560 30.240 91.820 ;
        RECT 30.340 91.560 30.600 91.820 ;
        RECT 30.700 91.560 30.960 91.820 ;
        RECT 31.060 91.560 31.320 91.820 ;
        RECT 31.420 91.560 31.680 91.820 ;
        RECT 31.780 91.560 32.040 91.820 ;
        RECT 32.140 91.560 32.400 91.820 ;
        RECT 32.500 91.560 32.760 91.820 ;
        RECT 32.860 91.560 33.120 91.820 ;
        RECT 33.220 91.560 33.480 91.820 ;
        RECT 33.580 91.560 33.840 91.820 ;
        RECT 33.940 91.560 34.200 91.820 ;
        RECT 34.300 91.560 34.560 91.820 ;
        RECT 34.660 91.560 34.920 91.820 ;
        RECT 35.020 91.560 35.280 91.820 ;
        RECT 35.380 91.560 35.640 91.820 ;
        RECT 35.740 91.560 36.000 91.820 ;
        RECT 36.100 91.560 36.360 91.820 ;
        RECT 36.460 91.560 36.720 91.820 ;
        RECT 36.820 91.560 37.080 91.820 ;
        RECT 37.180 91.560 37.440 91.820 ;
        RECT 37.540 91.560 37.800 91.820 ;
        RECT 37.900 91.560 38.160 91.820 ;
        RECT 38.260 91.560 38.520 91.820 ;
        RECT 38.620 91.560 38.880 91.820 ;
        RECT 38.980 91.560 39.240 91.820 ;
        RECT 39.340 91.560 39.600 91.820 ;
        RECT 39.700 91.560 39.960 91.820 ;
        RECT 40.060 91.560 40.320 91.820 ;
        RECT 40.420 91.560 40.680 91.820 ;
        RECT 40.780 91.560 41.040 91.820 ;
        RECT 41.140 91.560 41.400 91.820 ;
        RECT 41.500 91.560 41.760 91.820 ;
        RECT 41.860 91.560 42.120 91.820 ;
        RECT 42.220 91.560 42.480 91.820 ;
        RECT 42.580 91.560 42.840 91.820 ;
        RECT 42.940 91.560 43.200 91.820 ;
        RECT 43.300 91.560 43.560 91.820 ;
        RECT 43.660 91.560 43.920 91.820 ;
        RECT 44.020 91.560 44.280 91.820 ;
        RECT 44.380 91.560 44.640 91.820 ;
        RECT 44.740 91.560 45.000 91.820 ;
        RECT 45.100 91.560 45.360 91.820 ;
        RECT 45.460 91.560 45.720 91.820 ;
        RECT 45.820 91.560 46.080 91.820 ;
        RECT 46.180 91.560 46.440 91.820 ;
        RECT 46.540 91.560 46.800 91.820 ;
        RECT 46.900 91.560 47.160 91.820 ;
        RECT 47.260 91.560 47.520 91.820 ;
        RECT 47.620 91.560 47.880 91.820 ;
        RECT 47.980 91.560 48.240 91.820 ;
        RECT 48.340 91.560 48.600 91.820 ;
        RECT 48.700 91.560 48.960 91.820 ;
        RECT 49.060 91.560 49.320 91.820 ;
        RECT 49.420 91.560 49.680 91.820 ;
        RECT 49.780 91.560 50.040 91.820 ;
        RECT 50.140 91.560 50.400 91.820 ;
        RECT 50.500 91.560 50.760 91.820 ;
        RECT 50.860 91.560 51.120 91.820 ;
        RECT 51.220 91.560 51.480 91.820 ;
        RECT 11.620 91.200 11.880 91.460 ;
        RECT 11.980 91.200 12.240 91.460 ;
        RECT 12.340 91.200 12.600 91.460 ;
        RECT 12.700 91.200 12.960 91.460 ;
        RECT 13.060 91.200 13.320 91.460 ;
        RECT 13.420 91.200 13.680 91.460 ;
        RECT 13.780 91.200 14.040 91.460 ;
        RECT 14.140 91.200 14.400 91.460 ;
        RECT 14.500 91.200 14.760 91.460 ;
        RECT 14.860 91.200 15.120 91.460 ;
        RECT 15.220 91.200 15.480 91.460 ;
        RECT 15.580 91.200 15.840 91.460 ;
        RECT 15.940 91.200 16.200 91.460 ;
        RECT 16.300 91.200 16.560 91.460 ;
        RECT 16.660 91.200 16.920 91.460 ;
        RECT 17.020 91.200 17.280 91.460 ;
        RECT 17.380 91.200 17.640 91.460 ;
        RECT 17.740 91.200 18.000 91.460 ;
        RECT 18.100 91.200 18.360 91.460 ;
        RECT 18.460 91.200 18.720 91.460 ;
        RECT 18.820 91.200 19.080 91.460 ;
        RECT 19.180 91.200 19.440 91.460 ;
        RECT 19.540 91.200 19.800 91.460 ;
        RECT 19.900 91.200 20.160 91.460 ;
        RECT 20.260 91.200 20.520 91.460 ;
        RECT 20.620 91.200 20.880 91.460 ;
        RECT 20.980 91.200 21.240 91.460 ;
        RECT 21.340 91.200 21.600 91.460 ;
        RECT 21.700 91.200 21.960 91.460 ;
        RECT 22.060 91.200 22.320 91.460 ;
        RECT 22.420 91.200 22.680 91.460 ;
        RECT 22.780 91.200 23.040 91.460 ;
        RECT 23.140 91.200 23.400 91.460 ;
        RECT 23.500 91.200 23.760 91.460 ;
        RECT 23.860 91.200 24.120 91.460 ;
        RECT 24.220 91.200 24.480 91.460 ;
        RECT 24.580 91.200 24.840 91.460 ;
        RECT 24.940 91.200 25.200 91.460 ;
        RECT 25.300 91.200 25.560 91.460 ;
        RECT 25.660 91.200 25.920 91.460 ;
        RECT 26.020 91.200 26.280 91.460 ;
        RECT 26.380 91.200 26.640 91.460 ;
        RECT 26.740 91.200 27.000 91.460 ;
        RECT 27.100 91.200 27.360 91.460 ;
        RECT 27.460 91.200 27.720 91.460 ;
        RECT 27.820 91.200 28.080 91.460 ;
        RECT 28.180 91.200 28.440 91.460 ;
        RECT 28.540 91.200 28.800 91.460 ;
        RECT 28.900 91.200 29.160 91.460 ;
        RECT 29.260 91.200 29.520 91.460 ;
        RECT 29.620 91.200 29.880 91.460 ;
        RECT 29.980 91.200 30.240 91.460 ;
        RECT 30.340 91.200 30.600 91.460 ;
        RECT 30.700 91.200 30.960 91.460 ;
        RECT 31.060 91.200 31.320 91.460 ;
        RECT 31.420 91.200 31.680 91.460 ;
        RECT 31.780 91.200 32.040 91.460 ;
        RECT 32.140 91.200 32.400 91.460 ;
        RECT 32.500 91.200 32.760 91.460 ;
        RECT 32.860 91.200 33.120 91.460 ;
        RECT 33.220 91.200 33.480 91.460 ;
        RECT 33.580 91.200 33.840 91.460 ;
        RECT 33.940 91.200 34.200 91.460 ;
        RECT 34.300 91.200 34.560 91.460 ;
        RECT 34.660 91.200 34.920 91.460 ;
        RECT 35.020 91.200 35.280 91.460 ;
        RECT 35.380 91.200 35.640 91.460 ;
        RECT 35.740 91.200 36.000 91.460 ;
        RECT 36.100 91.200 36.360 91.460 ;
        RECT 36.460 91.200 36.720 91.460 ;
        RECT 36.820 91.200 37.080 91.460 ;
        RECT 37.180 91.200 37.440 91.460 ;
        RECT 37.540 91.200 37.800 91.460 ;
        RECT 37.900 91.200 38.160 91.460 ;
        RECT 38.260 91.200 38.520 91.460 ;
        RECT 38.620 91.200 38.880 91.460 ;
        RECT 38.980 91.200 39.240 91.460 ;
        RECT 39.340 91.200 39.600 91.460 ;
        RECT 39.700 91.200 39.960 91.460 ;
        RECT 40.060 91.200 40.320 91.460 ;
        RECT 40.420 91.200 40.680 91.460 ;
        RECT 40.780 91.200 41.040 91.460 ;
        RECT 41.140 91.200 41.400 91.460 ;
        RECT 41.500 91.200 41.760 91.460 ;
        RECT 41.860 91.200 42.120 91.460 ;
        RECT 42.220 91.200 42.480 91.460 ;
        RECT 42.580 91.200 42.840 91.460 ;
        RECT 42.940 91.200 43.200 91.460 ;
        RECT 43.300 91.200 43.560 91.460 ;
        RECT 43.660 91.200 43.920 91.460 ;
        RECT 44.020 91.200 44.280 91.460 ;
        RECT 44.380 91.200 44.640 91.460 ;
        RECT 44.740 91.200 45.000 91.460 ;
        RECT 45.100 91.200 45.360 91.460 ;
        RECT 45.460 91.200 45.720 91.460 ;
        RECT 45.820 91.200 46.080 91.460 ;
        RECT 46.180 91.200 46.440 91.460 ;
        RECT 46.540 91.200 46.800 91.460 ;
        RECT 46.900 91.200 47.160 91.460 ;
        RECT 47.260 91.200 47.520 91.460 ;
        RECT 47.620 91.200 47.880 91.460 ;
        RECT 47.980 91.200 48.240 91.460 ;
        RECT 48.340 91.200 48.600 91.460 ;
        RECT 48.700 91.200 48.960 91.460 ;
        RECT 49.060 91.200 49.320 91.460 ;
        RECT 49.420 91.200 49.680 91.460 ;
        RECT 49.780 91.200 50.040 91.460 ;
        RECT 50.140 91.200 50.400 91.460 ;
        RECT 50.500 91.200 50.760 91.460 ;
        RECT 50.860 91.200 51.120 91.460 ;
        RECT 51.220 91.200 51.480 91.460 ;
        RECT 11.620 90.840 11.880 91.100 ;
        RECT 11.980 90.840 12.240 91.100 ;
        RECT 12.340 90.840 12.600 91.100 ;
        RECT 12.700 90.840 12.960 91.100 ;
        RECT 13.060 90.840 13.320 91.100 ;
        RECT 13.420 90.840 13.680 91.100 ;
        RECT 13.780 90.840 14.040 91.100 ;
        RECT 14.140 90.840 14.400 91.100 ;
        RECT 14.500 90.840 14.760 91.100 ;
        RECT 14.860 90.840 15.120 91.100 ;
        RECT 15.220 90.840 15.480 91.100 ;
        RECT 15.580 90.840 15.840 91.100 ;
        RECT 15.940 90.840 16.200 91.100 ;
        RECT 16.300 90.840 16.560 91.100 ;
        RECT 16.660 90.840 16.920 91.100 ;
        RECT 17.020 90.840 17.280 91.100 ;
        RECT 17.380 90.840 17.640 91.100 ;
        RECT 17.740 90.840 18.000 91.100 ;
        RECT 18.100 90.840 18.360 91.100 ;
        RECT 18.460 90.840 18.720 91.100 ;
        RECT 18.820 90.840 19.080 91.100 ;
        RECT 19.180 90.840 19.440 91.100 ;
        RECT 19.540 90.840 19.800 91.100 ;
        RECT 19.900 90.840 20.160 91.100 ;
        RECT 20.260 90.840 20.520 91.100 ;
        RECT 20.620 90.840 20.880 91.100 ;
        RECT 20.980 90.840 21.240 91.100 ;
        RECT 21.340 90.840 21.600 91.100 ;
        RECT 21.700 90.840 21.960 91.100 ;
        RECT 22.060 90.840 22.320 91.100 ;
        RECT 22.420 90.840 22.680 91.100 ;
        RECT 22.780 90.840 23.040 91.100 ;
        RECT 23.140 90.840 23.400 91.100 ;
        RECT 23.500 90.840 23.760 91.100 ;
        RECT 23.860 90.840 24.120 91.100 ;
        RECT 24.220 90.840 24.480 91.100 ;
        RECT 24.580 90.840 24.840 91.100 ;
        RECT 24.940 90.840 25.200 91.100 ;
        RECT 25.300 90.840 25.560 91.100 ;
        RECT 25.660 90.840 25.920 91.100 ;
        RECT 26.020 90.840 26.280 91.100 ;
        RECT 26.380 90.840 26.640 91.100 ;
        RECT 26.740 90.840 27.000 91.100 ;
        RECT 27.100 90.840 27.360 91.100 ;
        RECT 27.460 90.840 27.720 91.100 ;
        RECT 27.820 90.840 28.080 91.100 ;
        RECT 28.180 90.840 28.440 91.100 ;
        RECT 28.540 90.840 28.800 91.100 ;
        RECT 28.900 90.840 29.160 91.100 ;
        RECT 29.260 90.840 29.520 91.100 ;
        RECT 29.620 90.840 29.880 91.100 ;
        RECT 29.980 90.840 30.240 91.100 ;
        RECT 30.340 90.840 30.600 91.100 ;
        RECT 30.700 90.840 30.960 91.100 ;
        RECT 31.060 90.840 31.320 91.100 ;
        RECT 31.420 90.840 31.680 91.100 ;
        RECT 31.780 90.840 32.040 91.100 ;
        RECT 32.140 90.840 32.400 91.100 ;
        RECT 32.500 90.840 32.760 91.100 ;
        RECT 32.860 90.840 33.120 91.100 ;
        RECT 33.220 90.840 33.480 91.100 ;
        RECT 33.580 90.840 33.840 91.100 ;
        RECT 33.940 90.840 34.200 91.100 ;
        RECT 34.300 90.840 34.560 91.100 ;
        RECT 34.660 90.840 34.920 91.100 ;
        RECT 35.020 90.840 35.280 91.100 ;
        RECT 35.380 90.840 35.640 91.100 ;
        RECT 35.740 90.840 36.000 91.100 ;
        RECT 36.100 90.840 36.360 91.100 ;
        RECT 36.460 90.840 36.720 91.100 ;
        RECT 36.820 90.840 37.080 91.100 ;
        RECT 37.180 90.840 37.440 91.100 ;
        RECT 37.540 90.840 37.800 91.100 ;
        RECT 37.900 90.840 38.160 91.100 ;
        RECT 38.260 90.840 38.520 91.100 ;
        RECT 38.620 90.840 38.880 91.100 ;
        RECT 38.980 90.840 39.240 91.100 ;
        RECT 39.340 90.840 39.600 91.100 ;
        RECT 39.700 90.840 39.960 91.100 ;
        RECT 40.060 90.840 40.320 91.100 ;
        RECT 40.420 90.840 40.680 91.100 ;
        RECT 40.780 90.840 41.040 91.100 ;
        RECT 41.140 90.840 41.400 91.100 ;
        RECT 41.500 90.840 41.760 91.100 ;
        RECT 41.860 90.840 42.120 91.100 ;
        RECT 42.220 90.840 42.480 91.100 ;
        RECT 42.580 90.840 42.840 91.100 ;
        RECT 42.940 90.840 43.200 91.100 ;
        RECT 43.300 90.840 43.560 91.100 ;
        RECT 43.660 90.840 43.920 91.100 ;
        RECT 44.020 90.840 44.280 91.100 ;
        RECT 44.380 90.840 44.640 91.100 ;
        RECT 44.740 90.840 45.000 91.100 ;
        RECT 45.100 90.840 45.360 91.100 ;
        RECT 45.460 90.840 45.720 91.100 ;
        RECT 45.820 90.840 46.080 91.100 ;
        RECT 46.180 90.840 46.440 91.100 ;
        RECT 46.540 90.840 46.800 91.100 ;
        RECT 46.900 90.840 47.160 91.100 ;
        RECT 47.260 90.840 47.520 91.100 ;
        RECT 47.620 90.840 47.880 91.100 ;
        RECT 47.980 90.840 48.240 91.100 ;
        RECT 48.340 90.840 48.600 91.100 ;
        RECT 48.700 90.840 48.960 91.100 ;
        RECT 49.060 90.840 49.320 91.100 ;
        RECT 49.420 90.840 49.680 91.100 ;
        RECT 49.780 90.840 50.040 91.100 ;
        RECT 50.140 90.840 50.400 91.100 ;
        RECT 50.500 90.840 50.760 91.100 ;
        RECT 50.860 90.840 51.120 91.100 ;
        RECT 51.220 90.840 51.480 91.100 ;
        RECT 56.850 89.660 57.110 89.920 ;
        RECT 57.210 89.660 57.470 89.920 ;
        RECT 57.570 89.660 57.830 89.920 ;
        RECT 57.930 89.660 58.190 89.920 ;
        RECT 58.290 89.660 58.550 89.920 ;
        RECT 58.650 89.660 58.910 89.920 ;
        RECT 59.010 89.660 59.270 89.920 ;
        RECT 59.370 89.660 59.630 89.920 ;
        RECT 59.730 89.660 59.990 89.920 ;
        RECT 60.090 89.660 60.350 89.920 ;
        RECT 60.450 89.660 60.710 89.920 ;
        RECT 60.810 89.660 61.070 89.920 ;
        RECT 61.170 89.660 61.430 89.920 ;
        RECT 61.530 89.660 61.790 89.920 ;
        RECT 61.890 89.660 62.150 89.920 ;
        RECT 62.250 89.660 62.510 89.920 ;
        RECT 62.610 89.660 62.870 89.920 ;
        RECT 62.970 89.660 63.230 89.920 ;
        RECT 63.330 89.660 63.590 89.920 ;
        RECT 63.690 89.660 63.950 89.920 ;
        RECT 64.050 89.660 64.310 89.920 ;
        RECT 64.410 89.660 64.670 89.920 ;
        RECT 64.770 89.660 65.030 89.920 ;
        RECT 65.130 89.660 65.390 89.920 ;
        RECT 65.490 89.660 65.750 89.920 ;
        RECT 65.850 89.660 66.110 89.920 ;
        RECT 66.210 89.660 66.470 89.920 ;
        RECT 66.570 89.660 66.830 89.920 ;
        RECT 66.930 89.660 67.190 89.920 ;
        RECT 67.290 89.660 67.550 89.920 ;
        RECT 67.650 89.660 67.910 89.920 ;
        RECT 68.010 89.660 68.270 89.920 ;
        RECT 68.370 89.660 68.630 89.920 ;
        RECT 68.730 89.660 68.990 89.920 ;
        RECT 69.090 89.660 69.350 89.920 ;
        RECT 69.450 89.660 69.710 89.920 ;
        RECT 69.810 89.660 70.070 89.920 ;
        RECT 70.170 89.660 70.430 89.920 ;
        RECT 70.530 89.660 70.790 89.920 ;
        RECT 70.890 89.660 71.150 89.920 ;
        RECT 71.250 89.660 71.510 89.920 ;
        RECT 71.610 89.660 71.870 89.920 ;
        RECT 71.970 89.660 72.230 89.920 ;
        RECT 72.330 89.660 72.590 89.920 ;
        RECT 72.690 89.660 72.950 89.920 ;
        RECT 73.050 89.660 73.310 89.920 ;
        RECT 73.410 89.660 73.670 89.920 ;
        RECT 73.770 89.660 74.030 89.920 ;
        RECT 74.130 89.660 74.390 89.920 ;
        RECT 74.490 89.660 74.750 89.920 ;
        RECT 74.850 89.660 75.110 89.920 ;
        RECT 75.210 89.660 75.470 89.920 ;
        RECT 75.570 89.660 75.830 89.920 ;
        RECT 75.930 89.660 76.190 89.920 ;
        RECT 76.290 89.660 76.550 89.920 ;
        RECT 76.650 89.660 76.910 89.920 ;
        RECT 77.010 89.660 77.270 89.920 ;
        RECT 77.370 89.660 77.630 89.920 ;
        RECT 77.730 89.660 77.990 89.920 ;
        RECT 78.090 89.660 78.350 89.920 ;
        RECT 78.450 89.660 78.710 89.920 ;
        RECT 78.810 89.660 79.070 89.920 ;
        RECT 79.170 89.660 79.430 89.920 ;
        RECT 79.530 89.660 79.790 89.920 ;
        RECT 79.890 89.660 80.150 89.920 ;
        RECT 80.250 89.660 80.510 89.920 ;
        RECT 80.610 89.660 80.870 89.920 ;
        RECT 80.970 89.660 81.230 89.920 ;
        RECT 81.330 89.660 81.590 89.920 ;
        RECT 81.690 89.660 81.950 89.920 ;
        RECT 82.050 89.660 82.310 89.920 ;
        RECT 82.410 89.660 82.670 89.920 ;
        RECT 82.770 89.660 83.030 89.920 ;
        RECT 83.130 89.660 83.390 89.920 ;
        RECT 83.490 89.660 83.750 89.920 ;
        RECT 83.850 89.660 84.110 89.920 ;
        RECT 84.210 89.660 84.470 89.920 ;
        RECT 84.570 89.660 84.830 89.920 ;
        RECT 84.930 89.660 85.190 89.920 ;
        RECT 85.290 89.660 85.550 89.920 ;
        RECT 85.650 89.660 85.910 89.920 ;
        RECT 86.010 89.660 86.270 89.920 ;
        RECT 86.370 89.660 86.630 89.920 ;
        RECT 86.730 89.660 86.990 89.920 ;
        RECT 87.090 89.660 87.350 89.920 ;
        RECT 87.450 89.660 87.710 89.920 ;
        RECT 87.810 89.660 88.070 89.920 ;
        RECT 88.170 89.660 88.430 89.920 ;
        RECT 88.530 89.660 88.790 89.920 ;
        RECT 88.890 89.660 89.150 89.920 ;
        RECT 89.250 89.660 89.510 89.920 ;
        RECT 89.610 89.660 89.870 89.920 ;
        RECT 89.970 89.660 90.230 89.920 ;
        RECT 90.330 89.660 90.590 89.920 ;
        RECT 90.690 89.660 90.950 89.920 ;
        RECT 91.050 89.660 91.310 89.920 ;
        RECT 91.410 89.660 91.670 89.920 ;
        RECT 91.770 89.660 92.030 89.920 ;
        RECT 92.130 89.660 92.390 89.920 ;
        RECT 92.490 89.660 92.750 89.920 ;
        RECT 92.850 89.660 93.110 89.920 ;
        RECT 93.210 89.660 93.470 89.920 ;
        RECT 93.570 89.660 93.830 89.920 ;
        RECT 93.930 89.660 94.190 89.920 ;
        RECT 94.290 89.660 94.550 89.920 ;
        RECT 94.650 89.660 94.910 89.920 ;
        RECT 95.010 89.660 95.270 89.920 ;
        RECT 95.370 89.660 95.630 89.920 ;
        RECT 95.730 89.660 95.990 89.920 ;
        RECT 96.090 89.660 96.350 89.920 ;
        RECT 96.450 89.660 96.710 89.920 ;
        RECT 56.850 89.300 57.110 89.560 ;
        RECT 57.210 89.300 57.470 89.560 ;
        RECT 57.570 89.300 57.830 89.560 ;
        RECT 57.930 89.300 58.190 89.560 ;
        RECT 58.290 89.300 58.550 89.560 ;
        RECT 58.650 89.300 58.910 89.560 ;
        RECT 59.010 89.300 59.270 89.560 ;
        RECT 59.370 89.300 59.630 89.560 ;
        RECT 59.730 89.300 59.990 89.560 ;
        RECT 60.090 89.300 60.350 89.560 ;
        RECT 60.450 89.300 60.710 89.560 ;
        RECT 60.810 89.300 61.070 89.560 ;
        RECT 61.170 89.300 61.430 89.560 ;
        RECT 61.530 89.300 61.790 89.560 ;
        RECT 61.890 89.300 62.150 89.560 ;
        RECT 62.250 89.300 62.510 89.560 ;
        RECT 62.610 89.300 62.870 89.560 ;
        RECT 62.970 89.300 63.230 89.560 ;
        RECT 63.330 89.300 63.590 89.560 ;
        RECT 63.690 89.300 63.950 89.560 ;
        RECT 64.050 89.300 64.310 89.560 ;
        RECT 64.410 89.300 64.670 89.560 ;
        RECT 64.770 89.300 65.030 89.560 ;
        RECT 65.130 89.300 65.390 89.560 ;
        RECT 65.490 89.300 65.750 89.560 ;
        RECT 65.850 89.300 66.110 89.560 ;
        RECT 66.210 89.300 66.470 89.560 ;
        RECT 66.570 89.300 66.830 89.560 ;
        RECT 66.930 89.300 67.190 89.560 ;
        RECT 67.290 89.300 67.550 89.560 ;
        RECT 67.650 89.300 67.910 89.560 ;
        RECT 68.010 89.300 68.270 89.560 ;
        RECT 68.370 89.300 68.630 89.560 ;
        RECT 68.730 89.300 68.990 89.560 ;
        RECT 69.090 89.300 69.350 89.560 ;
        RECT 69.450 89.300 69.710 89.560 ;
        RECT 69.810 89.300 70.070 89.560 ;
        RECT 70.170 89.300 70.430 89.560 ;
        RECT 70.530 89.300 70.790 89.560 ;
        RECT 70.890 89.300 71.150 89.560 ;
        RECT 71.250 89.300 71.510 89.560 ;
        RECT 71.610 89.300 71.870 89.560 ;
        RECT 71.970 89.300 72.230 89.560 ;
        RECT 72.330 89.300 72.590 89.560 ;
        RECT 72.690 89.300 72.950 89.560 ;
        RECT 73.050 89.300 73.310 89.560 ;
        RECT 73.410 89.300 73.670 89.560 ;
        RECT 73.770 89.300 74.030 89.560 ;
        RECT 74.130 89.300 74.390 89.560 ;
        RECT 74.490 89.300 74.750 89.560 ;
        RECT 74.850 89.300 75.110 89.560 ;
        RECT 75.210 89.300 75.470 89.560 ;
        RECT 75.570 89.300 75.830 89.560 ;
        RECT 75.930 89.300 76.190 89.560 ;
        RECT 76.290 89.300 76.550 89.560 ;
        RECT 76.650 89.300 76.910 89.560 ;
        RECT 77.010 89.300 77.270 89.560 ;
        RECT 77.370 89.300 77.630 89.560 ;
        RECT 77.730 89.300 77.990 89.560 ;
        RECT 78.090 89.300 78.350 89.560 ;
        RECT 78.450 89.300 78.710 89.560 ;
        RECT 78.810 89.300 79.070 89.560 ;
        RECT 79.170 89.300 79.430 89.560 ;
        RECT 79.530 89.300 79.790 89.560 ;
        RECT 79.890 89.300 80.150 89.560 ;
        RECT 80.250 89.300 80.510 89.560 ;
        RECT 80.610 89.300 80.870 89.560 ;
        RECT 80.970 89.300 81.230 89.560 ;
        RECT 81.330 89.300 81.590 89.560 ;
        RECT 81.690 89.300 81.950 89.560 ;
        RECT 82.050 89.300 82.310 89.560 ;
        RECT 82.410 89.300 82.670 89.560 ;
        RECT 82.770 89.300 83.030 89.560 ;
        RECT 83.130 89.300 83.390 89.560 ;
        RECT 83.490 89.300 83.750 89.560 ;
        RECT 83.850 89.300 84.110 89.560 ;
        RECT 84.210 89.300 84.470 89.560 ;
        RECT 84.570 89.300 84.830 89.560 ;
        RECT 84.930 89.300 85.190 89.560 ;
        RECT 85.290 89.300 85.550 89.560 ;
        RECT 85.650 89.300 85.910 89.560 ;
        RECT 86.010 89.300 86.270 89.560 ;
        RECT 86.370 89.300 86.630 89.560 ;
        RECT 86.730 89.300 86.990 89.560 ;
        RECT 87.090 89.300 87.350 89.560 ;
        RECT 87.450 89.300 87.710 89.560 ;
        RECT 87.810 89.300 88.070 89.560 ;
        RECT 88.170 89.300 88.430 89.560 ;
        RECT 88.530 89.300 88.790 89.560 ;
        RECT 88.890 89.300 89.150 89.560 ;
        RECT 89.250 89.300 89.510 89.560 ;
        RECT 89.610 89.300 89.870 89.560 ;
        RECT 89.970 89.300 90.230 89.560 ;
        RECT 90.330 89.300 90.590 89.560 ;
        RECT 90.690 89.300 90.950 89.560 ;
        RECT 91.050 89.300 91.310 89.560 ;
        RECT 91.410 89.300 91.670 89.560 ;
        RECT 91.770 89.300 92.030 89.560 ;
        RECT 92.130 89.300 92.390 89.560 ;
        RECT 92.490 89.300 92.750 89.560 ;
        RECT 92.850 89.300 93.110 89.560 ;
        RECT 93.210 89.300 93.470 89.560 ;
        RECT 93.570 89.300 93.830 89.560 ;
        RECT 93.930 89.300 94.190 89.560 ;
        RECT 94.290 89.300 94.550 89.560 ;
        RECT 94.650 89.300 94.910 89.560 ;
        RECT 95.010 89.300 95.270 89.560 ;
        RECT 95.370 89.300 95.630 89.560 ;
        RECT 95.730 89.300 95.990 89.560 ;
        RECT 96.090 89.300 96.350 89.560 ;
        RECT 96.450 89.300 96.710 89.560 ;
        RECT 56.850 88.940 57.110 89.200 ;
        RECT 57.210 88.940 57.470 89.200 ;
        RECT 57.570 88.940 57.830 89.200 ;
        RECT 57.930 88.940 58.190 89.200 ;
        RECT 58.290 88.940 58.550 89.200 ;
        RECT 58.650 88.940 58.910 89.200 ;
        RECT 59.010 88.940 59.270 89.200 ;
        RECT 59.370 88.940 59.630 89.200 ;
        RECT 59.730 88.940 59.990 89.200 ;
        RECT 60.090 88.940 60.350 89.200 ;
        RECT 60.450 88.940 60.710 89.200 ;
        RECT 60.810 88.940 61.070 89.200 ;
        RECT 61.170 88.940 61.430 89.200 ;
        RECT 61.530 88.940 61.790 89.200 ;
        RECT 61.890 88.940 62.150 89.200 ;
        RECT 62.250 88.940 62.510 89.200 ;
        RECT 62.610 88.940 62.870 89.200 ;
        RECT 62.970 88.940 63.230 89.200 ;
        RECT 63.330 88.940 63.590 89.200 ;
        RECT 63.690 88.940 63.950 89.200 ;
        RECT 64.050 88.940 64.310 89.200 ;
        RECT 64.410 88.940 64.670 89.200 ;
        RECT 64.770 88.940 65.030 89.200 ;
        RECT 65.130 88.940 65.390 89.200 ;
        RECT 65.490 88.940 65.750 89.200 ;
        RECT 65.850 88.940 66.110 89.200 ;
        RECT 66.210 88.940 66.470 89.200 ;
        RECT 66.570 88.940 66.830 89.200 ;
        RECT 66.930 88.940 67.190 89.200 ;
        RECT 67.290 88.940 67.550 89.200 ;
        RECT 67.650 88.940 67.910 89.200 ;
        RECT 68.010 88.940 68.270 89.200 ;
        RECT 68.370 88.940 68.630 89.200 ;
        RECT 68.730 88.940 68.990 89.200 ;
        RECT 69.090 88.940 69.350 89.200 ;
        RECT 69.450 88.940 69.710 89.200 ;
        RECT 69.810 88.940 70.070 89.200 ;
        RECT 70.170 88.940 70.430 89.200 ;
        RECT 70.530 88.940 70.790 89.200 ;
        RECT 70.890 88.940 71.150 89.200 ;
        RECT 71.250 88.940 71.510 89.200 ;
        RECT 71.610 88.940 71.870 89.200 ;
        RECT 71.970 88.940 72.230 89.200 ;
        RECT 72.330 88.940 72.590 89.200 ;
        RECT 72.690 88.940 72.950 89.200 ;
        RECT 73.050 88.940 73.310 89.200 ;
        RECT 73.410 88.940 73.670 89.200 ;
        RECT 73.770 88.940 74.030 89.200 ;
        RECT 74.130 88.940 74.390 89.200 ;
        RECT 74.490 88.940 74.750 89.200 ;
        RECT 74.850 88.940 75.110 89.200 ;
        RECT 75.210 88.940 75.470 89.200 ;
        RECT 75.570 88.940 75.830 89.200 ;
        RECT 75.930 88.940 76.190 89.200 ;
        RECT 76.290 88.940 76.550 89.200 ;
        RECT 76.650 88.940 76.910 89.200 ;
        RECT 77.010 88.940 77.270 89.200 ;
        RECT 77.370 88.940 77.630 89.200 ;
        RECT 77.730 88.940 77.990 89.200 ;
        RECT 78.090 88.940 78.350 89.200 ;
        RECT 78.450 88.940 78.710 89.200 ;
        RECT 78.810 88.940 79.070 89.200 ;
        RECT 79.170 88.940 79.430 89.200 ;
        RECT 79.530 88.940 79.790 89.200 ;
        RECT 79.890 88.940 80.150 89.200 ;
        RECT 80.250 88.940 80.510 89.200 ;
        RECT 80.610 88.940 80.870 89.200 ;
        RECT 80.970 88.940 81.230 89.200 ;
        RECT 81.330 88.940 81.590 89.200 ;
        RECT 81.690 88.940 81.950 89.200 ;
        RECT 82.050 88.940 82.310 89.200 ;
        RECT 82.410 88.940 82.670 89.200 ;
        RECT 82.770 88.940 83.030 89.200 ;
        RECT 83.130 88.940 83.390 89.200 ;
        RECT 83.490 88.940 83.750 89.200 ;
        RECT 83.850 88.940 84.110 89.200 ;
        RECT 84.210 88.940 84.470 89.200 ;
        RECT 84.570 88.940 84.830 89.200 ;
        RECT 84.930 88.940 85.190 89.200 ;
        RECT 85.290 88.940 85.550 89.200 ;
        RECT 85.650 88.940 85.910 89.200 ;
        RECT 86.010 88.940 86.270 89.200 ;
        RECT 86.370 88.940 86.630 89.200 ;
        RECT 86.730 88.940 86.990 89.200 ;
        RECT 87.090 88.940 87.350 89.200 ;
        RECT 87.450 88.940 87.710 89.200 ;
        RECT 87.810 88.940 88.070 89.200 ;
        RECT 88.170 88.940 88.430 89.200 ;
        RECT 88.530 88.940 88.790 89.200 ;
        RECT 88.890 88.940 89.150 89.200 ;
        RECT 89.250 88.940 89.510 89.200 ;
        RECT 89.610 88.940 89.870 89.200 ;
        RECT 89.970 88.940 90.230 89.200 ;
        RECT 90.330 88.940 90.590 89.200 ;
        RECT 90.690 88.940 90.950 89.200 ;
        RECT 91.050 88.940 91.310 89.200 ;
        RECT 91.410 88.940 91.670 89.200 ;
        RECT 91.770 88.940 92.030 89.200 ;
        RECT 92.130 88.940 92.390 89.200 ;
        RECT 92.490 88.940 92.750 89.200 ;
        RECT 92.850 88.940 93.110 89.200 ;
        RECT 93.210 88.940 93.470 89.200 ;
        RECT 93.570 88.940 93.830 89.200 ;
        RECT 93.930 88.940 94.190 89.200 ;
        RECT 94.290 88.940 94.550 89.200 ;
        RECT 94.650 88.940 94.910 89.200 ;
        RECT 95.010 88.940 95.270 89.200 ;
        RECT 95.370 88.940 95.630 89.200 ;
        RECT 95.730 88.940 95.990 89.200 ;
        RECT 96.090 88.940 96.350 89.200 ;
        RECT 96.450 88.940 96.710 89.200 ;
        RECT 100.335 88.950 100.595 89.210 ;
        RECT 100.695 88.950 100.955 89.210 ;
        RECT 101.055 88.950 101.315 89.210 ;
        RECT 100.335 88.590 100.595 88.850 ;
        RECT 100.695 88.590 100.955 88.850 ;
        RECT 101.055 88.590 101.315 88.850 ;
        RECT 100.335 88.230 100.595 88.490 ;
        RECT 100.695 88.230 100.955 88.490 ;
        RECT 101.055 88.230 101.315 88.490 ;
        RECT 16.530 87.585 16.790 87.845 ;
        RECT 16.890 87.585 17.150 87.845 ;
        RECT 17.250 87.585 17.510 87.845 ;
        RECT 16.530 87.225 16.790 87.485 ;
        RECT 16.890 87.225 17.150 87.485 ;
        RECT 17.250 87.225 17.510 87.485 ;
        RECT 16.530 86.865 16.790 87.125 ;
        RECT 16.890 86.865 17.150 87.125 ;
        RECT 17.250 86.865 17.510 87.125 ;
        RECT 16.530 86.505 16.790 86.765 ;
        RECT 16.890 86.505 17.150 86.765 ;
        RECT 17.250 86.505 17.510 86.765 ;
        RECT 16.530 86.145 16.790 86.405 ;
        RECT 16.890 86.145 17.150 86.405 ;
        RECT 17.250 86.145 17.510 86.405 ;
        RECT 16.530 85.785 16.790 86.045 ;
        RECT 16.890 85.785 17.150 86.045 ;
        RECT 17.250 85.785 17.510 86.045 ;
        RECT 16.530 85.425 16.790 85.685 ;
        RECT 16.890 85.425 17.150 85.685 ;
        RECT 17.250 85.425 17.510 85.685 ;
        RECT 16.530 85.065 16.790 85.325 ;
        RECT 16.890 85.065 17.150 85.325 ;
        RECT 17.250 85.065 17.510 85.325 ;
        RECT 16.530 84.705 16.790 84.965 ;
        RECT 16.890 84.705 17.150 84.965 ;
        RECT 17.250 84.705 17.510 84.965 ;
        RECT 16.530 84.345 16.790 84.605 ;
        RECT 16.890 84.345 17.150 84.605 ;
        RECT 17.250 84.345 17.510 84.605 ;
        RECT 16.530 83.985 16.790 84.245 ;
        RECT 16.890 83.985 17.150 84.245 ;
        RECT 17.250 83.985 17.510 84.245 ;
        RECT 16.530 83.625 16.790 83.885 ;
        RECT 16.890 83.625 17.150 83.885 ;
        RECT 17.250 83.625 17.510 83.885 ;
        RECT 16.530 83.265 16.790 83.525 ;
        RECT 16.890 83.265 17.150 83.525 ;
        RECT 17.250 83.265 17.510 83.525 ;
        RECT 16.530 82.905 16.790 83.165 ;
        RECT 16.890 82.905 17.150 83.165 ;
        RECT 17.250 82.905 17.510 83.165 ;
        RECT 16.530 82.545 16.790 82.805 ;
        RECT 16.890 82.545 17.150 82.805 ;
        RECT 17.250 82.545 17.510 82.805 ;
        RECT 16.530 82.185 16.790 82.445 ;
        RECT 16.890 82.185 17.150 82.445 ;
        RECT 17.250 82.185 17.510 82.445 ;
        RECT 16.530 81.825 16.790 82.085 ;
        RECT 16.890 81.825 17.150 82.085 ;
        RECT 17.250 81.825 17.510 82.085 ;
        RECT 16.530 81.465 16.790 81.725 ;
        RECT 16.890 81.465 17.150 81.725 ;
        RECT 17.250 81.465 17.510 81.725 ;
        RECT 16.530 81.105 16.790 81.365 ;
        RECT 16.890 81.105 17.150 81.365 ;
        RECT 17.250 81.105 17.510 81.365 ;
        RECT 16.530 80.745 16.790 81.005 ;
        RECT 16.890 80.745 17.150 81.005 ;
        RECT 17.250 80.745 17.510 81.005 ;
        RECT 16.530 80.385 16.790 80.645 ;
        RECT 16.890 80.385 17.150 80.645 ;
        RECT 17.250 80.385 17.510 80.645 ;
        RECT 16.530 80.025 16.790 80.285 ;
        RECT 16.890 80.025 17.150 80.285 ;
        RECT 17.250 80.025 17.510 80.285 ;
        RECT 16.530 79.665 16.790 79.925 ;
        RECT 16.890 79.665 17.150 79.925 ;
        RECT 17.250 79.665 17.510 79.925 ;
        RECT 16.530 79.305 16.790 79.565 ;
        RECT 16.890 79.305 17.150 79.565 ;
        RECT 17.250 79.305 17.510 79.565 ;
        RECT 16.530 78.945 16.790 79.205 ;
        RECT 16.890 78.945 17.150 79.205 ;
        RECT 17.250 78.945 17.510 79.205 ;
        RECT 16.530 78.585 16.790 78.845 ;
        RECT 16.890 78.585 17.150 78.845 ;
        RECT 17.250 78.585 17.510 78.845 ;
        RECT 16.530 78.225 16.790 78.485 ;
        RECT 16.890 78.225 17.150 78.485 ;
        RECT 17.250 78.225 17.510 78.485 ;
        RECT 16.530 77.865 16.790 78.125 ;
        RECT 16.890 77.865 17.150 78.125 ;
        RECT 17.250 77.865 17.510 78.125 ;
        RECT 16.530 77.505 16.790 77.765 ;
        RECT 16.890 77.505 17.150 77.765 ;
        RECT 17.250 77.505 17.510 77.765 ;
        RECT 16.530 77.145 16.790 77.405 ;
        RECT 16.890 77.145 17.150 77.405 ;
        RECT 17.250 77.145 17.510 77.405 ;
        RECT 16.530 76.785 16.790 77.045 ;
        RECT 16.890 76.785 17.150 77.045 ;
        RECT 17.250 76.785 17.510 77.045 ;
        RECT 16.530 76.425 16.790 76.685 ;
        RECT 16.890 76.425 17.150 76.685 ;
        RECT 17.250 76.425 17.510 76.685 ;
        RECT 16.530 76.065 16.790 76.325 ;
        RECT 16.890 76.065 17.150 76.325 ;
        RECT 17.250 76.065 17.510 76.325 ;
        RECT 16.530 75.705 16.790 75.965 ;
        RECT 16.890 75.705 17.150 75.965 ;
        RECT 17.250 75.705 17.510 75.965 ;
        RECT 16.530 75.345 16.790 75.605 ;
        RECT 16.890 75.345 17.150 75.605 ;
        RECT 17.250 75.345 17.510 75.605 ;
        RECT 16.530 74.985 16.790 75.245 ;
        RECT 16.890 74.985 17.150 75.245 ;
        RECT 17.250 74.985 17.510 75.245 ;
        RECT 16.530 74.625 16.790 74.885 ;
        RECT 16.890 74.625 17.150 74.885 ;
        RECT 17.250 74.625 17.510 74.885 ;
        RECT 16.530 74.265 16.790 74.525 ;
        RECT 16.890 74.265 17.150 74.525 ;
        RECT 17.250 74.265 17.510 74.525 ;
        RECT 16.530 73.905 16.790 74.165 ;
        RECT 16.890 73.905 17.150 74.165 ;
        RECT 17.250 73.905 17.510 74.165 ;
        RECT 16.530 73.545 16.790 73.805 ;
        RECT 16.890 73.545 17.150 73.805 ;
        RECT 17.250 73.545 17.510 73.805 ;
        RECT 16.530 73.185 16.790 73.445 ;
        RECT 16.890 73.185 17.150 73.445 ;
        RECT 17.250 73.185 17.510 73.445 ;
        RECT 16.530 72.825 16.790 73.085 ;
        RECT 16.890 72.825 17.150 73.085 ;
        RECT 17.250 72.825 17.510 73.085 ;
        RECT 16.530 72.465 16.790 72.725 ;
        RECT 16.890 72.465 17.150 72.725 ;
        RECT 17.250 72.465 17.510 72.725 ;
        RECT 16.530 72.105 16.790 72.365 ;
        RECT 16.890 72.105 17.150 72.365 ;
        RECT 17.250 72.105 17.510 72.365 ;
        RECT 16.530 71.745 16.790 72.005 ;
        RECT 16.890 71.745 17.150 72.005 ;
        RECT 17.250 71.745 17.510 72.005 ;
        RECT 16.530 71.385 16.790 71.645 ;
        RECT 16.890 71.385 17.150 71.645 ;
        RECT 17.250 71.385 17.510 71.645 ;
        RECT 16.530 71.025 16.790 71.285 ;
        RECT 16.890 71.025 17.150 71.285 ;
        RECT 17.250 71.025 17.510 71.285 ;
        RECT 16.530 70.665 16.790 70.925 ;
        RECT 16.890 70.665 17.150 70.925 ;
        RECT 17.250 70.665 17.510 70.925 ;
        RECT 16.530 70.305 16.790 70.565 ;
        RECT 16.890 70.305 17.150 70.565 ;
        RECT 17.250 70.305 17.510 70.565 ;
        RECT 16.530 69.945 16.790 70.205 ;
        RECT 16.890 69.945 17.150 70.205 ;
        RECT 17.250 69.945 17.510 70.205 ;
        RECT 16.530 69.585 16.790 69.845 ;
        RECT 16.890 69.585 17.150 69.845 ;
        RECT 17.250 69.585 17.510 69.845 ;
        RECT 16.530 69.225 16.790 69.485 ;
        RECT 16.890 69.225 17.150 69.485 ;
        RECT 17.250 69.225 17.510 69.485 ;
        RECT 16.530 68.865 16.790 69.125 ;
        RECT 16.890 68.865 17.150 69.125 ;
        RECT 17.250 68.865 17.510 69.125 ;
        RECT 16.530 68.505 16.790 68.765 ;
        RECT 16.890 68.505 17.150 68.765 ;
        RECT 17.250 68.505 17.510 68.765 ;
        RECT 16.530 68.145 16.790 68.405 ;
        RECT 16.890 68.145 17.150 68.405 ;
        RECT 17.250 68.145 17.510 68.405 ;
        RECT 16.530 67.785 16.790 68.045 ;
        RECT 16.890 67.785 17.150 68.045 ;
        RECT 17.250 67.785 17.510 68.045 ;
        RECT 16.530 67.425 16.790 67.685 ;
        RECT 16.890 67.425 17.150 67.685 ;
        RECT 17.250 67.425 17.510 67.685 ;
        RECT 16.530 67.065 16.790 67.325 ;
        RECT 16.890 67.065 17.150 67.325 ;
        RECT 17.250 67.065 17.510 67.325 ;
        RECT 16.530 66.705 16.790 66.965 ;
        RECT 16.890 66.705 17.150 66.965 ;
        RECT 17.250 66.705 17.510 66.965 ;
        RECT 16.530 66.345 16.790 66.605 ;
        RECT 16.890 66.345 17.150 66.605 ;
        RECT 17.250 66.345 17.510 66.605 ;
        RECT 16.530 65.985 16.790 66.245 ;
        RECT 16.890 65.985 17.150 66.245 ;
        RECT 17.250 65.985 17.510 66.245 ;
        RECT 16.530 65.625 16.790 65.885 ;
        RECT 16.890 65.625 17.150 65.885 ;
        RECT 17.250 65.625 17.510 65.885 ;
        RECT 16.530 65.265 16.790 65.525 ;
        RECT 16.890 65.265 17.150 65.525 ;
        RECT 17.250 65.265 17.510 65.525 ;
        RECT 16.530 64.905 16.790 65.165 ;
        RECT 16.890 64.905 17.150 65.165 ;
        RECT 17.250 64.905 17.510 65.165 ;
        RECT 16.530 64.545 16.790 64.805 ;
        RECT 16.890 64.545 17.150 64.805 ;
        RECT 17.250 64.545 17.510 64.805 ;
        RECT 16.530 64.185 16.790 64.445 ;
        RECT 16.890 64.185 17.150 64.445 ;
        RECT 17.250 64.185 17.510 64.445 ;
        RECT 16.530 63.825 16.790 64.085 ;
        RECT 16.890 63.825 17.150 64.085 ;
        RECT 17.250 63.825 17.510 64.085 ;
        RECT 16.530 63.465 16.790 63.725 ;
        RECT 16.890 63.465 17.150 63.725 ;
        RECT 17.250 63.465 17.510 63.725 ;
        RECT 16.530 63.105 16.790 63.365 ;
        RECT 16.890 63.105 17.150 63.365 ;
        RECT 17.250 63.105 17.510 63.365 ;
        RECT 16.530 62.745 16.790 63.005 ;
        RECT 16.890 62.745 17.150 63.005 ;
        RECT 17.250 62.745 17.510 63.005 ;
        RECT 16.530 62.385 16.790 62.645 ;
        RECT 16.890 62.385 17.150 62.645 ;
        RECT 17.250 62.385 17.510 62.645 ;
        RECT 16.530 62.025 16.790 62.285 ;
        RECT 16.890 62.025 17.150 62.285 ;
        RECT 17.250 62.025 17.510 62.285 ;
        RECT 16.530 61.665 16.790 61.925 ;
        RECT 16.890 61.665 17.150 61.925 ;
        RECT 17.250 61.665 17.510 61.925 ;
        RECT 16.530 61.305 16.790 61.565 ;
        RECT 16.890 61.305 17.150 61.565 ;
        RECT 17.250 61.305 17.510 61.565 ;
        RECT 16.530 60.945 16.790 61.205 ;
        RECT 16.890 60.945 17.150 61.205 ;
        RECT 17.250 60.945 17.510 61.205 ;
        RECT 16.530 60.585 16.790 60.845 ;
        RECT 16.890 60.585 17.150 60.845 ;
        RECT 17.250 60.585 17.510 60.845 ;
        RECT 16.530 60.225 16.790 60.485 ;
        RECT 16.890 60.225 17.150 60.485 ;
        RECT 17.250 60.225 17.510 60.485 ;
        RECT 16.530 59.865 16.790 60.125 ;
        RECT 16.890 59.865 17.150 60.125 ;
        RECT 17.250 59.865 17.510 60.125 ;
        RECT 16.530 59.505 16.790 59.765 ;
        RECT 16.890 59.505 17.150 59.765 ;
        RECT 17.250 59.505 17.510 59.765 ;
        RECT 16.530 59.145 16.790 59.405 ;
        RECT 16.890 59.145 17.150 59.405 ;
        RECT 17.250 59.145 17.510 59.405 ;
        RECT 16.530 58.785 16.790 59.045 ;
        RECT 16.890 58.785 17.150 59.045 ;
        RECT 17.250 58.785 17.510 59.045 ;
        RECT 16.530 58.425 16.790 58.685 ;
        RECT 16.890 58.425 17.150 58.685 ;
        RECT 17.250 58.425 17.510 58.685 ;
        RECT 16.530 58.065 16.790 58.325 ;
        RECT 16.890 58.065 17.150 58.325 ;
        RECT 17.250 58.065 17.510 58.325 ;
        RECT 16.530 57.705 16.790 57.965 ;
        RECT 16.890 57.705 17.150 57.965 ;
        RECT 17.250 57.705 17.510 57.965 ;
        RECT 16.530 57.345 16.790 57.605 ;
        RECT 16.890 57.345 17.150 57.605 ;
        RECT 17.250 57.345 17.510 57.605 ;
        RECT 16.530 56.985 16.790 57.245 ;
        RECT 16.890 56.985 17.150 57.245 ;
        RECT 17.250 56.985 17.510 57.245 ;
        RECT 16.530 56.625 16.790 56.885 ;
        RECT 16.890 56.625 17.150 56.885 ;
        RECT 17.250 56.625 17.510 56.885 ;
        RECT 16.530 56.265 16.790 56.525 ;
        RECT 16.890 56.265 17.150 56.525 ;
        RECT 17.250 56.265 17.510 56.525 ;
        RECT 16.530 55.905 16.790 56.165 ;
        RECT 16.890 55.905 17.150 56.165 ;
        RECT 17.250 55.905 17.510 56.165 ;
        RECT 16.530 55.545 16.790 55.805 ;
        RECT 16.890 55.545 17.150 55.805 ;
        RECT 17.250 55.545 17.510 55.805 ;
        RECT 16.530 55.185 16.790 55.445 ;
        RECT 16.890 55.185 17.150 55.445 ;
        RECT 17.250 55.185 17.510 55.445 ;
        RECT 16.530 54.825 16.790 55.085 ;
        RECT 16.890 54.825 17.150 55.085 ;
        RECT 17.250 54.825 17.510 55.085 ;
        RECT 16.530 54.465 16.790 54.725 ;
        RECT 16.890 54.465 17.150 54.725 ;
        RECT 17.250 54.465 17.510 54.725 ;
        RECT 16.530 54.105 16.790 54.365 ;
        RECT 16.890 54.105 17.150 54.365 ;
        RECT 17.250 54.105 17.510 54.365 ;
        RECT 16.530 53.745 16.790 54.005 ;
        RECT 16.890 53.745 17.150 54.005 ;
        RECT 17.250 53.745 17.510 54.005 ;
        RECT 16.530 53.385 16.790 53.645 ;
        RECT 16.890 53.385 17.150 53.645 ;
        RECT 17.250 53.385 17.510 53.645 ;
        RECT 16.530 53.025 16.790 53.285 ;
        RECT 16.890 53.025 17.150 53.285 ;
        RECT 17.250 53.025 17.510 53.285 ;
        RECT 16.530 52.665 16.790 52.925 ;
        RECT 16.890 52.665 17.150 52.925 ;
        RECT 17.250 52.665 17.510 52.925 ;
        RECT 16.530 52.305 16.790 52.565 ;
        RECT 16.890 52.305 17.150 52.565 ;
        RECT 17.250 52.305 17.510 52.565 ;
        RECT 16.530 51.945 16.790 52.205 ;
        RECT 16.890 51.945 17.150 52.205 ;
        RECT 17.250 51.945 17.510 52.205 ;
        RECT 16.530 51.585 16.790 51.845 ;
        RECT 16.890 51.585 17.150 51.845 ;
        RECT 17.250 51.585 17.510 51.845 ;
        RECT 16.530 51.225 16.790 51.485 ;
        RECT 16.890 51.225 17.150 51.485 ;
        RECT 17.250 51.225 17.510 51.485 ;
        RECT 16.530 50.865 16.790 51.125 ;
        RECT 16.890 50.865 17.150 51.125 ;
        RECT 17.250 50.865 17.510 51.125 ;
        RECT 16.530 50.505 16.790 50.765 ;
        RECT 16.890 50.505 17.150 50.765 ;
        RECT 17.250 50.505 17.510 50.765 ;
        RECT 16.530 50.145 16.790 50.405 ;
        RECT 16.890 50.145 17.150 50.405 ;
        RECT 17.250 50.145 17.510 50.405 ;
        RECT 16.530 49.785 16.790 50.045 ;
        RECT 16.890 49.785 17.150 50.045 ;
        RECT 17.250 49.785 17.510 50.045 ;
        RECT 16.530 49.425 16.790 49.685 ;
        RECT 16.890 49.425 17.150 49.685 ;
        RECT 17.250 49.425 17.510 49.685 ;
        RECT 16.530 49.065 16.790 49.325 ;
        RECT 16.890 49.065 17.150 49.325 ;
        RECT 17.250 49.065 17.510 49.325 ;
        RECT 100.335 87.870 100.595 88.130 ;
        RECT 100.695 87.870 100.955 88.130 ;
        RECT 101.055 87.870 101.315 88.130 ;
        RECT 100.335 87.510 100.595 87.770 ;
        RECT 100.695 87.510 100.955 87.770 ;
        RECT 101.055 87.510 101.315 87.770 ;
        RECT 100.335 87.150 100.595 87.410 ;
        RECT 100.695 87.150 100.955 87.410 ;
        RECT 101.055 87.150 101.315 87.410 ;
        RECT 100.335 86.790 100.595 87.050 ;
        RECT 100.695 86.790 100.955 87.050 ;
        RECT 101.055 86.790 101.315 87.050 ;
        RECT 100.335 86.430 100.595 86.690 ;
        RECT 100.695 86.430 100.955 86.690 ;
        RECT 101.055 86.430 101.315 86.690 ;
        RECT 100.335 86.070 100.595 86.330 ;
        RECT 100.695 86.070 100.955 86.330 ;
        RECT 101.055 86.070 101.315 86.330 ;
        RECT 100.335 85.710 100.595 85.970 ;
        RECT 100.695 85.710 100.955 85.970 ;
        RECT 101.055 85.710 101.315 85.970 ;
        RECT 100.335 85.350 100.595 85.610 ;
        RECT 100.695 85.350 100.955 85.610 ;
        RECT 101.055 85.350 101.315 85.610 ;
        RECT 100.335 84.990 100.595 85.250 ;
        RECT 100.695 84.990 100.955 85.250 ;
        RECT 101.055 84.990 101.315 85.250 ;
        RECT 100.335 84.630 100.595 84.890 ;
        RECT 100.695 84.630 100.955 84.890 ;
        RECT 101.055 84.630 101.315 84.890 ;
        RECT 100.335 84.270 100.595 84.530 ;
        RECT 100.695 84.270 100.955 84.530 ;
        RECT 101.055 84.270 101.315 84.530 ;
        RECT 100.335 83.910 100.595 84.170 ;
        RECT 100.695 83.910 100.955 84.170 ;
        RECT 101.055 83.910 101.315 84.170 ;
        RECT 100.335 83.550 100.595 83.810 ;
        RECT 100.695 83.550 100.955 83.810 ;
        RECT 101.055 83.550 101.315 83.810 ;
        RECT 100.335 83.190 100.595 83.450 ;
        RECT 100.695 83.190 100.955 83.450 ;
        RECT 101.055 83.190 101.315 83.450 ;
        RECT 100.335 82.830 100.595 83.090 ;
        RECT 100.695 82.830 100.955 83.090 ;
        RECT 101.055 82.830 101.315 83.090 ;
        RECT 100.335 82.470 100.595 82.730 ;
        RECT 100.695 82.470 100.955 82.730 ;
        RECT 101.055 82.470 101.315 82.730 ;
        RECT 100.335 82.110 100.595 82.370 ;
        RECT 100.695 82.110 100.955 82.370 ;
        RECT 101.055 82.110 101.315 82.370 ;
        RECT 100.335 81.750 100.595 82.010 ;
        RECT 100.695 81.750 100.955 82.010 ;
        RECT 101.055 81.750 101.315 82.010 ;
        RECT 100.335 81.390 100.595 81.650 ;
        RECT 100.695 81.390 100.955 81.650 ;
        RECT 101.055 81.390 101.315 81.650 ;
        RECT 100.335 81.030 100.595 81.290 ;
        RECT 100.695 81.030 100.955 81.290 ;
        RECT 101.055 81.030 101.315 81.290 ;
        RECT 100.335 80.670 100.595 80.930 ;
        RECT 100.695 80.670 100.955 80.930 ;
        RECT 101.055 80.670 101.315 80.930 ;
        RECT 100.335 80.310 100.595 80.570 ;
        RECT 100.695 80.310 100.955 80.570 ;
        RECT 101.055 80.310 101.315 80.570 ;
        RECT 100.335 79.950 100.595 80.210 ;
        RECT 100.695 79.950 100.955 80.210 ;
        RECT 101.055 79.950 101.315 80.210 ;
        RECT 100.335 79.590 100.595 79.850 ;
        RECT 100.695 79.590 100.955 79.850 ;
        RECT 101.055 79.590 101.315 79.850 ;
        RECT 100.335 79.230 100.595 79.490 ;
        RECT 100.695 79.230 100.955 79.490 ;
        RECT 101.055 79.230 101.315 79.490 ;
        RECT 100.335 78.870 100.595 79.130 ;
        RECT 100.695 78.870 100.955 79.130 ;
        RECT 101.055 78.870 101.315 79.130 ;
        RECT 100.335 78.510 100.595 78.770 ;
        RECT 100.695 78.510 100.955 78.770 ;
        RECT 101.055 78.510 101.315 78.770 ;
        RECT 100.335 78.150 100.595 78.410 ;
        RECT 100.695 78.150 100.955 78.410 ;
        RECT 101.055 78.150 101.315 78.410 ;
        RECT 100.335 77.790 100.595 78.050 ;
        RECT 100.695 77.790 100.955 78.050 ;
        RECT 101.055 77.790 101.315 78.050 ;
        RECT 100.335 77.430 100.595 77.690 ;
        RECT 100.695 77.430 100.955 77.690 ;
        RECT 101.055 77.430 101.315 77.690 ;
        RECT 100.335 77.070 100.595 77.330 ;
        RECT 100.695 77.070 100.955 77.330 ;
        RECT 101.055 77.070 101.315 77.330 ;
        RECT 100.335 76.710 100.595 76.970 ;
        RECT 100.695 76.710 100.955 76.970 ;
        RECT 101.055 76.710 101.315 76.970 ;
        RECT 100.335 76.350 100.595 76.610 ;
        RECT 100.695 76.350 100.955 76.610 ;
        RECT 101.055 76.350 101.315 76.610 ;
        RECT 100.335 75.990 100.595 76.250 ;
        RECT 100.695 75.990 100.955 76.250 ;
        RECT 101.055 75.990 101.315 76.250 ;
        RECT 100.335 75.630 100.595 75.890 ;
        RECT 100.695 75.630 100.955 75.890 ;
        RECT 101.055 75.630 101.315 75.890 ;
        RECT 100.335 75.270 100.595 75.530 ;
        RECT 100.695 75.270 100.955 75.530 ;
        RECT 101.055 75.270 101.315 75.530 ;
        RECT 100.335 74.910 100.595 75.170 ;
        RECT 100.695 74.910 100.955 75.170 ;
        RECT 101.055 74.910 101.315 75.170 ;
        RECT 100.335 74.550 100.595 74.810 ;
        RECT 100.695 74.550 100.955 74.810 ;
        RECT 101.055 74.550 101.315 74.810 ;
        RECT 100.335 74.190 100.595 74.450 ;
        RECT 100.695 74.190 100.955 74.450 ;
        RECT 101.055 74.190 101.315 74.450 ;
        RECT 100.335 73.830 100.595 74.090 ;
        RECT 100.695 73.830 100.955 74.090 ;
        RECT 101.055 73.830 101.315 74.090 ;
        RECT 100.335 73.470 100.595 73.730 ;
        RECT 100.695 73.470 100.955 73.730 ;
        RECT 101.055 73.470 101.315 73.730 ;
        RECT 100.335 73.110 100.595 73.370 ;
        RECT 100.695 73.110 100.955 73.370 ;
        RECT 101.055 73.110 101.315 73.370 ;
        RECT 100.335 72.750 100.595 73.010 ;
        RECT 100.695 72.750 100.955 73.010 ;
        RECT 101.055 72.750 101.315 73.010 ;
        RECT 100.335 72.390 100.595 72.650 ;
        RECT 100.695 72.390 100.955 72.650 ;
        RECT 101.055 72.390 101.315 72.650 ;
        RECT 100.335 72.030 100.595 72.290 ;
        RECT 100.695 72.030 100.955 72.290 ;
        RECT 101.055 72.030 101.315 72.290 ;
        RECT 100.335 71.670 100.595 71.930 ;
        RECT 100.695 71.670 100.955 71.930 ;
        RECT 101.055 71.670 101.315 71.930 ;
        RECT 100.335 71.310 100.595 71.570 ;
        RECT 100.695 71.310 100.955 71.570 ;
        RECT 101.055 71.310 101.315 71.570 ;
        RECT 100.335 70.950 100.595 71.210 ;
        RECT 100.695 70.950 100.955 71.210 ;
        RECT 101.055 70.950 101.315 71.210 ;
        RECT 100.335 70.590 100.595 70.850 ;
        RECT 100.695 70.590 100.955 70.850 ;
        RECT 101.055 70.590 101.315 70.850 ;
        RECT 100.335 70.230 100.595 70.490 ;
        RECT 100.695 70.230 100.955 70.490 ;
        RECT 101.055 70.230 101.315 70.490 ;
        RECT 100.335 69.870 100.595 70.130 ;
        RECT 100.695 69.870 100.955 70.130 ;
        RECT 101.055 69.870 101.315 70.130 ;
        RECT 100.335 69.510 100.595 69.770 ;
        RECT 100.695 69.510 100.955 69.770 ;
        RECT 101.055 69.510 101.315 69.770 ;
        RECT 100.335 69.150 100.595 69.410 ;
        RECT 100.695 69.150 100.955 69.410 ;
        RECT 101.055 69.150 101.315 69.410 ;
        RECT 100.335 68.790 100.595 69.050 ;
        RECT 100.695 68.790 100.955 69.050 ;
        RECT 101.055 68.790 101.315 69.050 ;
        RECT 100.335 68.430 100.595 68.690 ;
        RECT 100.695 68.430 100.955 68.690 ;
        RECT 101.055 68.430 101.315 68.690 ;
        RECT 100.335 68.070 100.595 68.330 ;
        RECT 100.695 68.070 100.955 68.330 ;
        RECT 101.055 68.070 101.315 68.330 ;
        RECT 100.335 67.710 100.595 67.970 ;
        RECT 100.695 67.710 100.955 67.970 ;
        RECT 101.055 67.710 101.315 67.970 ;
        RECT 100.335 67.350 100.595 67.610 ;
        RECT 100.695 67.350 100.955 67.610 ;
        RECT 101.055 67.350 101.315 67.610 ;
        RECT 100.335 66.990 100.595 67.250 ;
        RECT 100.695 66.990 100.955 67.250 ;
        RECT 101.055 66.990 101.315 67.250 ;
        RECT 100.335 66.630 100.595 66.890 ;
        RECT 100.695 66.630 100.955 66.890 ;
        RECT 101.055 66.630 101.315 66.890 ;
        RECT 100.335 66.270 100.595 66.530 ;
        RECT 100.695 66.270 100.955 66.530 ;
        RECT 101.055 66.270 101.315 66.530 ;
        RECT 100.335 65.910 100.595 66.170 ;
        RECT 100.695 65.910 100.955 66.170 ;
        RECT 101.055 65.910 101.315 66.170 ;
        RECT 100.335 65.550 100.595 65.810 ;
        RECT 100.695 65.550 100.955 65.810 ;
        RECT 101.055 65.550 101.315 65.810 ;
        RECT 100.335 65.190 100.595 65.450 ;
        RECT 100.695 65.190 100.955 65.450 ;
        RECT 101.055 65.190 101.315 65.450 ;
        RECT 100.335 64.830 100.595 65.090 ;
        RECT 100.695 64.830 100.955 65.090 ;
        RECT 101.055 64.830 101.315 65.090 ;
        RECT 100.335 64.470 100.595 64.730 ;
        RECT 100.695 64.470 100.955 64.730 ;
        RECT 101.055 64.470 101.315 64.730 ;
        RECT 100.335 64.110 100.595 64.370 ;
        RECT 100.695 64.110 100.955 64.370 ;
        RECT 101.055 64.110 101.315 64.370 ;
        RECT 100.335 63.750 100.595 64.010 ;
        RECT 100.695 63.750 100.955 64.010 ;
        RECT 101.055 63.750 101.315 64.010 ;
        RECT 100.335 63.390 100.595 63.650 ;
        RECT 100.695 63.390 100.955 63.650 ;
        RECT 101.055 63.390 101.315 63.650 ;
        RECT 100.335 63.030 100.595 63.290 ;
        RECT 100.695 63.030 100.955 63.290 ;
        RECT 101.055 63.030 101.315 63.290 ;
        RECT 100.335 62.670 100.595 62.930 ;
        RECT 100.695 62.670 100.955 62.930 ;
        RECT 101.055 62.670 101.315 62.930 ;
        RECT 100.335 62.310 100.595 62.570 ;
        RECT 100.695 62.310 100.955 62.570 ;
        RECT 101.055 62.310 101.315 62.570 ;
        RECT 100.335 61.950 100.595 62.210 ;
        RECT 100.695 61.950 100.955 62.210 ;
        RECT 101.055 61.950 101.315 62.210 ;
        RECT 100.335 61.590 100.595 61.850 ;
        RECT 100.695 61.590 100.955 61.850 ;
        RECT 101.055 61.590 101.315 61.850 ;
        RECT 100.335 61.230 100.595 61.490 ;
        RECT 100.695 61.230 100.955 61.490 ;
        RECT 101.055 61.230 101.315 61.490 ;
        RECT 100.335 60.870 100.595 61.130 ;
        RECT 100.695 60.870 100.955 61.130 ;
        RECT 101.055 60.870 101.315 61.130 ;
        RECT 100.335 60.510 100.595 60.770 ;
        RECT 100.695 60.510 100.955 60.770 ;
        RECT 101.055 60.510 101.315 60.770 ;
        RECT 100.335 60.150 100.595 60.410 ;
        RECT 100.695 60.150 100.955 60.410 ;
        RECT 101.055 60.150 101.315 60.410 ;
        RECT 100.335 59.790 100.595 60.050 ;
        RECT 100.695 59.790 100.955 60.050 ;
        RECT 101.055 59.790 101.315 60.050 ;
        RECT 100.335 59.430 100.595 59.690 ;
        RECT 100.695 59.430 100.955 59.690 ;
        RECT 101.055 59.430 101.315 59.690 ;
        RECT 100.335 59.070 100.595 59.330 ;
        RECT 100.695 59.070 100.955 59.330 ;
        RECT 101.055 59.070 101.315 59.330 ;
        RECT 100.335 58.710 100.595 58.970 ;
        RECT 100.695 58.710 100.955 58.970 ;
        RECT 101.055 58.710 101.315 58.970 ;
        RECT 100.335 58.350 100.595 58.610 ;
        RECT 100.695 58.350 100.955 58.610 ;
        RECT 101.055 58.350 101.315 58.610 ;
        RECT 100.335 57.990 100.595 58.250 ;
        RECT 100.695 57.990 100.955 58.250 ;
        RECT 101.055 57.990 101.315 58.250 ;
        RECT 100.335 57.630 100.595 57.890 ;
        RECT 100.695 57.630 100.955 57.890 ;
        RECT 101.055 57.630 101.315 57.890 ;
        RECT 100.335 57.270 100.595 57.530 ;
        RECT 100.695 57.270 100.955 57.530 ;
        RECT 101.055 57.270 101.315 57.530 ;
        RECT 100.335 56.910 100.595 57.170 ;
        RECT 100.695 56.910 100.955 57.170 ;
        RECT 101.055 56.910 101.315 57.170 ;
        RECT 100.335 56.550 100.595 56.810 ;
        RECT 100.695 56.550 100.955 56.810 ;
        RECT 101.055 56.550 101.315 56.810 ;
        RECT 100.335 56.190 100.595 56.450 ;
        RECT 100.695 56.190 100.955 56.450 ;
        RECT 101.055 56.190 101.315 56.450 ;
        RECT 100.335 55.830 100.595 56.090 ;
        RECT 100.695 55.830 100.955 56.090 ;
        RECT 101.055 55.830 101.315 56.090 ;
        RECT 100.335 55.470 100.595 55.730 ;
        RECT 100.695 55.470 100.955 55.730 ;
        RECT 101.055 55.470 101.315 55.730 ;
        RECT 100.335 55.110 100.595 55.370 ;
        RECT 100.695 55.110 100.955 55.370 ;
        RECT 101.055 55.110 101.315 55.370 ;
        RECT 100.335 54.750 100.595 55.010 ;
        RECT 100.695 54.750 100.955 55.010 ;
        RECT 101.055 54.750 101.315 55.010 ;
        RECT 100.335 54.390 100.595 54.650 ;
        RECT 100.695 54.390 100.955 54.650 ;
        RECT 101.055 54.390 101.315 54.650 ;
        RECT 100.335 54.030 100.595 54.290 ;
        RECT 100.695 54.030 100.955 54.290 ;
        RECT 101.055 54.030 101.315 54.290 ;
        RECT 100.335 53.670 100.595 53.930 ;
        RECT 100.695 53.670 100.955 53.930 ;
        RECT 101.055 53.670 101.315 53.930 ;
        RECT 100.335 53.310 100.595 53.570 ;
        RECT 100.695 53.310 100.955 53.570 ;
        RECT 101.055 53.310 101.315 53.570 ;
        RECT 100.335 52.950 100.595 53.210 ;
        RECT 100.695 52.950 100.955 53.210 ;
        RECT 101.055 52.950 101.315 53.210 ;
        RECT 100.335 52.590 100.595 52.850 ;
        RECT 100.695 52.590 100.955 52.850 ;
        RECT 101.055 52.590 101.315 52.850 ;
        RECT 100.335 52.230 100.595 52.490 ;
        RECT 100.695 52.230 100.955 52.490 ;
        RECT 101.055 52.230 101.315 52.490 ;
        RECT 100.335 51.870 100.595 52.130 ;
        RECT 100.695 51.870 100.955 52.130 ;
        RECT 101.055 51.870 101.315 52.130 ;
        RECT 100.335 51.510 100.595 51.770 ;
        RECT 100.695 51.510 100.955 51.770 ;
        RECT 101.055 51.510 101.315 51.770 ;
        RECT 100.335 51.150 100.595 51.410 ;
        RECT 100.695 51.150 100.955 51.410 ;
        RECT 101.055 51.150 101.315 51.410 ;
        RECT 100.335 50.790 100.595 51.050 ;
        RECT 100.695 50.790 100.955 51.050 ;
        RECT 101.055 50.790 101.315 51.050 ;
        RECT 100.335 50.430 100.595 50.690 ;
        RECT 100.695 50.430 100.955 50.690 ;
        RECT 101.055 50.430 101.315 50.690 ;
        RECT 100.335 50.070 100.595 50.330 ;
        RECT 100.695 50.070 100.955 50.330 ;
        RECT 101.055 50.070 101.315 50.330 ;
        RECT 100.335 49.710 100.595 49.970 ;
        RECT 100.695 49.710 100.955 49.970 ;
        RECT 101.055 49.710 101.315 49.970 ;
        RECT 100.335 49.350 100.595 49.610 ;
        RECT 100.695 49.350 100.955 49.610 ;
        RECT 101.055 49.350 101.315 49.610 ;
        RECT 16.530 48.705 16.790 48.965 ;
        RECT 16.890 48.705 17.150 48.965 ;
        RECT 17.250 48.705 17.510 48.965 ;
        RECT 16.530 48.345 16.790 48.605 ;
        RECT 16.890 48.345 17.150 48.605 ;
        RECT 17.250 48.345 17.510 48.605 ;
        RECT 16.530 47.985 16.790 48.245 ;
        RECT 16.890 47.985 17.150 48.245 ;
        RECT 17.250 47.985 17.510 48.245 ;
        RECT 22.580 45.330 22.840 45.590 ;
        RECT 22.940 45.330 23.200 45.590 ;
        RECT 23.300 45.330 23.560 45.590 ;
        RECT 22.580 44.970 22.840 45.230 ;
        RECT 22.940 44.970 23.200 45.230 ;
        RECT 23.300 44.970 23.560 45.230 ;
        RECT 22.580 44.610 22.840 44.870 ;
        RECT 22.940 44.610 23.200 44.870 ;
        RECT 23.300 44.610 23.560 44.870 ;
        RECT 22.580 44.250 22.840 44.510 ;
        RECT 22.940 44.250 23.200 44.510 ;
        RECT 23.300 44.250 23.560 44.510 ;
        RECT 22.580 43.890 22.840 44.150 ;
        RECT 22.940 43.890 23.200 44.150 ;
        RECT 23.300 43.890 23.560 44.150 ;
        RECT 22.580 43.530 22.840 43.790 ;
        RECT 22.940 43.530 23.200 43.790 ;
        RECT 23.300 43.530 23.560 43.790 ;
        RECT 22.580 43.170 22.840 43.430 ;
        RECT 22.940 43.170 23.200 43.430 ;
        RECT 23.300 43.170 23.560 43.430 ;
        RECT 22.580 42.810 22.840 43.070 ;
        RECT 22.940 42.810 23.200 43.070 ;
        RECT 23.300 42.810 23.560 43.070 ;
        RECT 22.580 42.450 22.840 42.710 ;
        RECT 22.940 42.450 23.200 42.710 ;
        RECT 23.300 42.450 23.560 42.710 ;
        RECT 22.580 42.090 22.840 42.350 ;
        RECT 22.940 42.090 23.200 42.350 ;
        RECT 23.300 42.090 23.560 42.350 ;
        RECT 22.580 41.730 22.840 41.990 ;
        RECT 22.940 41.730 23.200 41.990 ;
        RECT 23.300 41.730 23.560 41.990 ;
        RECT 22.580 41.370 22.840 41.630 ;
        RECT 22.940 41.370 23.200 41.630 ;
        RECT 23.300 41.370 23.560 41.630 ;
        RECT 22.580 41.010 22.840 41.270 ;
        RECT 22.940 41.010 23.200 41.270 ;
        RECT 23.300 41.010 23.560 41.270 ;
        RECT 22.580 40.650 22.840 40.910 ;
        RECT 22.940 40.650 23.200 40.910 ;
        RECT 23.300 40.650 23.560 40.910 ;
        RECT 22.580 40.290 22.840 40.550 ;
        RECT 22.940 40.290 23.200 40.550 ;
        RECT 23.300 40.290 23.560 40.550 ;
        RECT 22.580 39.930 22.840 40.190 ;
        RECT 22.940 39.930 23.200 40.190 ;
        RECT 23.300 39.930 23.560 40.190 ;
        RECT 22.580 39.570 22.840 39.830 ;
        RECT 22.940 39.570 23.200 39.830 ;
        RECT 23.300 39.570 23.560 39.830 ;
        RECT 22.580 39.210 22.840 39.470 ;
        RECT 22.940 39.210 23.200 39.470 ;
        RECT 23.300 39.210 23.560 39.470 ;
        RECT 22.580 38.850 22.840 39.110 ;
        RECT 22.940 38.850 23.200 39.110 ;
        RECT 23.300 38.850 23.560 39.110 ;
        RECT 22.580 38.490 22.840 38.750 ;
        RECT 22.940 38.490 23.200 38.750 ;
        RECT 23.300 38.490 23.560 38.750 ;
        RECT 22.580 38.130 22.840 38.390 ;
        RECT 22.940 38.130 23.200 38.390 ;
        RECT 23.300 38.130 23.560 38.390 ;
        RECT 22.580 37.770 22.840 38.030 ;
        RECT 22.940 37.770 23.200 38.030 ;
        RECT 23.300 37.770 23.560 38.030 ;
        RECT 22.580 37.410 22.840 37.670 ;
        RECT 22.940 37.410 23.200 37.670 ;
        RECT 23.300 37.410 23.560 37.670 ;
        RECT 22.580 37.050 22.840 37.310 ;
        RECT 22.940 37.050 23.200 37.310 ;
        RECT 23.300 37.050 23.560 37.310 ;
        RECT 22.580 36.690 22.840 36.950 ;
        RECT 22.940 36.690 23.200 36.950 ;
        RECT 23.300 36.690 23.560 36.950 ;
        RECT 22.580 36.330 22.840 36.590 ;
        RECT 22.940 36.330 23.200 36.590 ;
        RECT 23.300 36.330 23.560 36.590 ;
        RECT 22.580 35.970 22.840 36.230 ;
        RECT 22.940 35.970 23.200 36.230 ;
        RECT 23.300 35.970 23.560 36.230 ;
        RECT 22.580 35.610 22.840 35.870 ;
        RECT 22.940 35.610 23.200 35.870 ;
        RECT 23.300 35.610 23.560 35.870 ;
        RECT 22.580 35.250 22.840 35.510 ;
        RECT 22.940 35.250 23.200 35.510 ;
        RECT 23.300 35.250 23.560 35.510 ;
        RECT 22.580 34.890 22.840 35.150 ;
        RECT 22.940 34.890 23.200 35.150 ;
        RECT 23.300 34.890 23.560 35.150 ;
        RECT 22.580 34.530 22.840 34.790 ;
        RECT 22.940 34.530 23.200 34.790 ;
        RECT 23.300 34.530 23.560 34.790 ;
        RECT 22.580 34.170 22.840 34.430 ;
        RECT 22.940 34.170 23.200 34.430 ;
        RECT 23.300 34.170 23.560 34.430 ;
        RECT 22.580 33.810 22.840 34.070 ;
        RECT 22.940 33.810 23.200 34.070 ;
        RECT 23.300 33.810 23.560 34.070 ;
        RECT 22.580 33.450 22.840 33.710 ;
        RECT 22.940 33.450 23.200 33.710 ;
        RECT 23.300 33.450 23.560 33.710 ;
        RECT 22.580 33.090 22.840 33.350 ;
        RECT 22.940 33.090 23.200 33.350 ;
        RECT 23.300 33.090 23.560 33.350 ;
        RECT 22.580 32.730 22.840 32.990 ;
        RECT 22.940 32.730 23.200 32.990 ;
        RECT 23.300 32.730 23.560 32.990 ;
        RECT 22.580 32.370 22.840 32.630 ;
        RECT 22.940 32.370 23.200 32.630 ;
        RECT 23.300 32.370 23.560 32.630 ;
        RECT 22.580 32.010 22.840 32.270 ;
        RECT 22.940 32.010 23.200 32.270 ;
        RECT 23.300 32.010 23.560 32.270 ;
        RECT 22.580 31.650 22.840 31.910 ;
        RECT 22.940 31.650 23.200 31.910 ;
        RECT 23.300 31.650 23.560 31.910 ;
        RECT 22.580 31.290 22.840 31.550 ;
        RECT 22.940 31.290 23.200 31.550 ;
        RECT 23.300 31.290 23.560 31.550 ;
        RECT 22.580 30.930 22.840 31.190 ;
        RECT 22.940 30.930 23.200 31.190 ;
        RECT 23.300 30.930 23.560 31.190 ;
        RECT 22.580 30.570 22.840 30.830 ;
        RECT 22.940 30.570 23.200 30.830 ;
        RECT 23.300 30.570 23.560 30.830 ;
        RECT 22.580 30.210 22.840 30.470 ;
        RECT 22.940 30.210 23.200 30.470 ;
        RECT 23.300 30.210 23.560 30.470 ;
        RECT 22.580 29.850 22.840 30.110 ;
        RECT 22.940 29.850 23.200 30.110 ;
        RECT 23.300 29.850 23.560 30.110 ;
        RECT 22.580 29.490 22.840 29.750 ;
        RECT 22.940 29.490 23.200 29.750 ;
        RECT 23.300 29.490 23.560 29.750 ;
        RECT 22.580 29.130 22.840 29.390 ;
        RECT 22.940 29.130 23.200 29.390 ;
        RECT 23.300 29.130 23.560 29.390 ;
        RECT 22.580 28.770 22.840 29.030 ;
        RECT 22.940 28.770 23.200 29.030 ;
        RECT 23.300 28.770 23.560 29.030 ;
        RECT 22.580 28.410 22.840 28.670 ;
        RECT 22.940 28.410 23.200 28.670 ;
        RECT 23.300 28.410 23.560 28.670 ;
        RECT 22.580 28.050 22.840 28.310 ;
        RECT 22.940 28.050 23.200 28.310 ;
        RECT 23.300 28.050 23.560 28.310 ;
        RECT 22.580 27.690 22.840 27.950 ;
        RECT 22.940 27.690 23.200 27.950 ;
        RECT 23.300 27.690 23.560 27.950 ;
        RECT 22.580 27.330 22.840 27.590 ;
        RECT 22.940 27.330 23.200 27.590 ;
        RECT 23.300 27.330 23.560 27.590 ;
        RECT 22.580 26.970 22.840 27.230 ;
        RECT 22.940 26.970 23.200 27.230 ;
        RECT 23.300 26.970 23.560 27.230 ;
        RECT 66.365 27.605 66.625 27.865 ;
        RECT 66.725 27.605 66.985 27.865 ;
        RECT 67.085 27.605 67.345 27.865 ;
        RECT 67.445 27.605 67.705 27.865 ;
        RECT 67.805 27.605 68.065 27.865 ;
        RECT 68.165 27.605 68.425 27.865 ;
        RECT 68.525 27.605 68.785 27.865 ;
        RECT 68.885 27.605 69.145 27.865 ;
        RECT 69.245 27.605 69.505 27.865 ;
        RECT 69.605 27.605 69.865 27.865 ;
        RECT 69.965 27.605 70.225 27.865 ;
        RECT 70.325 27.605 70.585 27.865 ;
        RECT 70.685 27.605 70.945 27.865 ;
        RECT 71.045 27.605 71.305 27.865 ;
        RECT 71.405 27.605 71.665 27.865 ;
        RECT 71.765 27.605 72.025 27.865 ;
        RECT 72.125 27.605 72.385 27.865 ;
        RECT 72.485 27.605 72.745 27.865 ;
        RECT 72.845 27.605 73.105 27.865 ;
        RECT 73.205 27.605 73.465 27.865 ;
        RECT 73.565 27.605 73.825 27.865 ;
        RECT 73.925 27.605 74.185 27.865 ;
        RECT 74.285 27.605 74.545 27.865 ;
        RECT 74.645 27.605 74.905 27.865 ;
        RECT 75.005 27.605 75.265 27.865 ;
        RECT 75.365 27.605 75.625 27.865 ;
        RECT 75.725 27.605 75.985 27.865 ;
        RECT 76.085 27.605 76.345 27.865 ;
        RECT 76.445 27.605 76.705 27.865 ;
        RECT 76.805 27.605 77.065 27.865 ;
        RECT 77.165 27.605 77.425 27.865 ;
        RECT 77.525 27.605 77.785 27.865 ;
        RECT 77.885 27.605 78.145 27.865 ;
        RECT 78.245 27.605 78.505 27.865 ;
        RECT 78.605 27.605 78.865 27.865 ;
        RECT 78.965 27.605 79.225 27.865 ;
        RECT 79.325 27.605 79.585 27.865 ;
        RECT 79.685 27.605 79.945 27.865 ;
        RECT 80.045 27.605 80.305 27.865 ;
        RECT 80.405 27.605 80.665 27.865 ;
        RECT 80.765 27.605 81.025 27.865 ;
        RECT 81.125 27.605 81.385 27.865 ;
        RECT 81.485 27.605 81.745 27.865 ;
        RECT 81.845 27.605 82.105 27.865 ;
        RECT 82.205 27.605 82.465 27.865 ;
        RECT 82.565 27.605 82.825 27.865 ;
        RECT 82.925 27.605 83.185 27.865 ;
        RECT 83.285 27.605 83.545 27.865 ;
        RECT 83.645 27.605 83.905 27.865 ;
        RECT 84.005 27.605 84.265 27.865 ;
        RECT 84.365 27.605 84.625 27.865 ;
        RECT 84.725 27.605 84.985 27.865 ;
        RECT 85.085 27.605 85.345 27.865 ;
        RECT 85.445 27.605 85.705 27.865 ;
        RECT 85.805 27.605 86.065 27.865 ;
        RECT 86.165 27.605 86.425 27.865 ;
        RECT 86.525 27.605 86.785 27.865 ;
        RECT 86.885 27.605 87.145 27.865 ;
        RECT 87.245 27.605 87.505 27.865 ;
        RECT 87.605 27.605 87.865 27.865 ;
        RECT 87.965 27.605 88.225 27.865 ;
        RECT 88.325 27.605 88.585 27.865 ;
        RECT 88.685 27.605 88.945 27.865 ;
        RECT 89.045 27.605 89.305 27.865 ;
        RECT 89.405 27.605 89.665 27.865 ;
        RECT 89.765 27.605 90.025 27.865 ;
        RECT 90.125 27.605 90.385 27.865 ;
        RECT 90.485 27.605 90.745 27.865 ;
        RECT 90.845 27.605 91.105 27.865 ;
        RECT 91.205 27.605 91.465 27.865 ;
        RECT 91.565 27.605 91.825 27.865 ;
        RECT 91.925 27.605 92.185 27.865 ;
        RECT 92.285 27.605 92.545 27.865 ;
        RECT 92.645 27.605 92.905 27.865 ;
        RECT 93.005 27.605 93.265 27.865 ;
        RECT 93.365 27.605 93.625 27.865 ;
        RECT 93.725 27.605 93.985 27.865 ;
        RECT 94.085 27.605 94.345 27.865 ;
        RECT 94.445 27.605 94.705 27.865 ;
        RECT 94.805 27.605 95.065 27.865 ;
        RECT 95.165 27.605 95.425 27.865 ;
        RECT 95.525 27.605 95.785 27.865 ;
        RECT 95.885 27.605 96.145 27.865 ;
        RECT 96.245 27.605 96.505 27.865 ;
        RECT 96.605 27.605 96.865 27.865 ;
        RECT 96.965 27.605 97.225 27.865 ;
        RECT 97.325 27.605 97.585 27.865 ;
        RECT 97.685 27.605 97.945 27.865 ;
        RECT 98.045 27.605 98.305 27.865 ;
        RECT 98.405 27.605 98.665 27.865 ;
        RECT 98.765 27.605 99.025 27.865 ;
        RECT 99.125 27.605 99.385 27.865 ;
        RECT 99.485 27.605 99.745 27.865 ;
        RECT 99.845 27.605 100.105 27.865 ;
        RECT 100.205 27.605 100.465 27.865 ;
        RECT 100.565 27.605 100.825 27.865 ;
        RECT 100.925 27.605 101.185 27.865 ;
        RECT 101.285 27.605 101.545 27.865 ;
        RECT 101.645 27.605 101.905 27.865 ;
        RECT 102.005 27.605 102.265 27.865 ;
        RECT 102.365 27.605 102.625 27.865 ;
        RECT 102.725 27.605 102.985 27.865 ;
        RECT 103.085 27.605 103.345 27.865 ;
        RECT 103.445 27.605 103.705 27.865 ;
        RECT 103.805 27.605 104.065 27.865 ;
        RECT 104.165 27.605 104.425 27.865 ;
        RECT 104.525 27.605 104.785 27.865 ;
        RECT 104.885 27.605 105.145 27.865 ;
        RECT 105.245 27.605 105.505 27.865 ;
        RECT 105.605 27.605 105.865 27.865 ;
        RECT 105.965 27.605 106.225 27.865 ;
        RECT 66.365 27.245 66.625 27.505 ;
        RECT 66.725 27.245 66.985 27.505 ;
        RECT 67.085 27.245 67.345 27.505 ;
        RECT 67.445 27.245 67.705 27.505 ;
        RECT 67.805 27.245 68.065 27.505 ;
        RECT 68.165 27.245 68.425 27.505 ;
        RECT 68.525 27.245 68.785 27.505 ;
        RECT 68.885 27.245 69.145 27.505 ;
        RECT 69.245 27.245 69.505 27.505 ;
        RECT 69.605 27.245 69.865 27.505 ;
        RECT 69.965 27.245 70.225 27.505 ;
        RECT 70.325 27.245 70.585 27.505 ;
        RECT 70.685 27.245 70.945 27.505 ;
        RECT 71.045 27.245 71.305 27.505 ;
        RECT 71.405 27.245 71.665 27.505 ;
        RECT 71.765 27.245 72.025 27.505 ;
        RECT 72.125 27.245 72.385 27.505 ;
        RECT 72.485 27.245 72.745 27.505 ;
        RECT 72.845 27.245 73.105 27.505 ;
        RECT 73.205 27.245 73.465 27.505 ;
        RECT 73.565 27.245 73.825 27.505 ;
        RECT 73.925 27.245 74.185 27.505 ;
        RECT 74.285 27.245 74.545 27.505 ;
        RECT 74.645 27.245 74.905 27.505 ;
        RECT 75.005 27.245 75.265 27.505 ;
        RECT 75.365 27.245 75.625 27.505 ;
        RECT 75.725 27.245 75.985 27.505 ;
        RECT 76.085 27.245 76.345 27.505 ;
        RECT 76.445 27.245 76.705 27.505 ;
        RECT 76.805 27.245 77.065 27.505 ;
        RECT 77.165 27.245 77.425 27.505 ;
        RECT 77.525 27.245 77.785 27.505 ;
        RECT 77.885 27.245 78.145 27.505 ;
        RECT 78.245 27.245 78.505 27.505 ;
        RECT 78.605 27.245 78.865 27.505 ;
        RECT 78.965 27.245 79.225 27.505 ;
        RECT 79.325 27.245 79.585 27.505 ;
        RECT 79.685 27.245 79.945 27.505 ;
        RECT 80.045 27.245 80.305 27.505 ;
        RECT 80.405 27.245 80.665 27.505 ;
        RECT 80.765 27.245 81.025 27.505 ;
        RECT 81.125 27.245 81.385 27.505 ;
        RECT 81.485 27.245 81.745 27.505 ;
        RECT 81.845 27.245 82.105 27.505 ;
        RECT 82.205 27.245 82.465 27.505 ;
        RECT 82.565 27.245 82.825 27.505 ;
        RECT 82.925 27.245 83.185 27.505 ;
        RECT 83.285 27.245 83.545 27.505 ;
        RECT 83.645 27.245 83.905 27.505 ;
        RECT 84.005 27.245 84.265 27.505 ;
        RECT 84.365 27.245 84.625 27.505 ;
        RECT 84.725 27.245 84.985 27.505 ;
        RECT 85.085 27.245 85.345 27.505 ;
        RECT 85.445 27.245 85.705 27.505 ;
        RECT 85.805 27.245 86.065 27.505 ;
        RECT 86.165 27.245 86.425 27.505 ;
        RECT 86.525 27.245 86.785 27.505 ;
        RECT 86.885 27.245 87.145 27.505 ;
        RECT 87.245 27.245 87.505 27.505 ;
        RECT 87.605 27.245 87.865 27.505 ;
        RECT 87.965 27.245 88.225 27.505 ;
        RECT 88.325 27.245 88.585 27.505 ;
        RECT 88.685 27.245 88.945 27.505 ;
        RECT 89.045 27.245 89.305 27.505 ;
        RECT 89.405 27.245 89.665 27.505 ;
        RECT 89.765 27.245 90.025 27.505 ;
        RECT 90.125 27.245 90.385 27.505 ;
        RECT 90.485 27.245 90.745 27.505 ;
        RECT 90.845 27.245 91.105 27.505 ;
        RECT 91.205 27.245 91.465 27.505 ;
        RECT 91.565 27.245 91.825 27.505 ;
        RECT 91.925 27.245 92.185 27.505 ;
        RECT 92.285 27.245 92.545 27.505 ;
        RECT 92.645 27.245 92.905 27.505 ;
        RECT 93.005 27.245 93.265 27.505 ;
        RECT 93.365 27.245 93.625 27.505 ;
        RECT 93.725 27.245 93.985 27.505 ;
        RECT 94.085 27.245 94.345 27.505 ;
        RECT 94.445 27.245 94.705 27.505 ;
        RECT 94.805 27.245 95.065 27.505 ;
        RECT 95.165 27.245 95.425 27.505 ;
        RECT 95.525 27.245 95.785 27.505 ;
        RECT 95.885 27.245 96.145 27.505 ;
        RECT 96.245 27.245 96.505 27.505 ;
        RECT 96.605 27.245 96.865 27.505 ;
        RECT 96.965 27.245 97.225 27.505 ;
        RECT 97.325 27.245 97.585 27.505 ;
        RECT 97.685 27.245 97.945 27.505 ;
        RECT 98.045 27.245 98.305 27.505 ;
        RECT 98.405 27.245 98.665 27.505 ;
        RECT 98.765 27.245 99.025 27.505 ;
        RECT 99.125 27.245 99.385 27.505 ;
        RECT 99.485 27.245 99.745 27.505 ;
        RECT 99.845 27.245 100.105 27.505 ;
        RECT 100.205 27.245 100.465 27.505 ;
        RECT 100.565 27.245 100.825 27.505 ;
        RECT 100.925 27.245 101.185 27.505 ;
        RECT 101.285 27.245 101.545 27.505 ;
        RECT 101.645 27.245 101.905 27.505 ;
        RECT 102.005 27.245 102.265 27.505 ;
        RECT 102.365 27.245 102.625 27.505 ;
        RECT 102.725 27.245 102.985 27.505 ;
        RECT 103.085 27.245 103.345 27.505 ;
        RECT 103.445 27.245 103.705 27.505 ;
        RECT 103.805 27.245 104.065 27.505 ;
        RECT 104.165 27.245 104.425 27.505 ;
        RECT 104.525 27.245 104.785 27.505 ;
        RECT 104.885 27.245 105.145 27.505 ;
        RECT 105.245 27.245 105.505 27.505 ;
        RECT 105.605 27.245 105.865 27.505 ;
        RECT 105.965 27.245 106.225 27.505 ;
        RECT 22.580 26.610 22.840 26.870 ;
        RECT 22.940 26.610 23.200 26.870 ;
        RECT 23.300 26.610 23.560 26.870 ;
        RECT 22.580 26.250 22.840 26.510 ;
        RECT 22.940 26.250 23.200 26.510 ;
        RECT 23.300 26.250 23.560 26.510 ;
        RECT 22.580 25.890 22.840 26.150 ;
        RECT 22.940 25.890 23.200 26.150 ;
        RECT 23.300 25.890 23.560 26.150 ;
        RECT 22.580 25.530 22.840 25.790 ;
        RECT 22.940 25.530 23.200 25.790 ;
        RECT 23.300 25.530 23.560 25.790 ;
        RECT 66.365 26.885 66.625 27.145 ;
        RECT 66.725 26.885 66.985 27.145 ;
        RECT 67.085 26.885 67.345 27.145 ;
        RECT 67.445 26.885 67.705 27.145 ;
        RECT 67.805 26.885 68.065 27.145 ;
        RECT 68.165 26.885 68.425 27.145 ;
        RECT 68.525 26.885 68.785 27.145 ;
        RECT 68.885 26.885 69.145 27.145 ;
        RECT 69.245 26.885 69.505 27.145 ;
        RECT 69.605 26.885 69.865 27.145 ;
        RECT 69.965 26.885 70.225 27.145 ;
        RECT 70.325 26.885 70.585 27.145 ;
        RECT 70.685 26.885 70.945 27.145 ;
        RECT 71.045 26.885 71.305 27.145 ;
        RECT 71.405 26.885 71.665 27.145 ;
        RECT 71.765 26.885 72.025 27.145 ;
        RECT 72.125 26.885 72.385 27.145 ;
        RECT 72.485 26.885 72.745 27.145 ;
        RECT 72.845 26.885 73.105 27.145 ;
        RECT 73.205 26.885 73.465 27.145 ;
        RECT 73.565 26.885 73.825 27.145 ;
        RECT 73.925 26.885 74.185 27.145 ;
        RECT 74.285 26.885 74.545 27.145 ;
        RECT 74.645 26.885 74.905 27.145 ;
        RECT 75.005 26.885 75.265 27.145 ;
        RECT 75.365 26.885 75.625 27.145 ;
        RECT 75.725 26.885 75.985 27.145 ;
        RECT 76.085 26.885 76.345 27.145 ;
        RECT 76.445 26.885 76.705 27.145 ;
        RECT 76.805 26.885 77.065 27.145 ;
        RECT 77.165 26.885 77.425 27.145 ;
        RECT 77.525 26.885 77.785 27.145 ;
        RECT 77.885 26.885 78.145 27.145 ;
        RECT 78.245 26.885 78.505 27.145 ;
        RECT 78.605 26.885 78.865 27.145 ;
        RECT 78.965 26.885 79.225 27.145 ;
        RECT 79.325 26.885 79.585 27.145 ;
        RECT 79.685 26.885 79.945 27.145 ;
        RECT 80.045 26.885 80.305 27.145 ;
        RECT 80.405 26.885 80.665 27.145 ;
        RECT 80.765 26.885 81.025 27.145 ;
        RECT 81.125 26.885 81.385 27.145 ;
        RECT 81.485 26.885 81.745 27.145 ;
        RECT 81.845 26.885 82.105 27.145 ;
        RECT 82.205 26.885 82.465 27.145 ;
        RECT 82.565 26.885 82.825 27.145 ;
        RECT 82.925 26.885 83.185 27.145 ;
        RECT 83.285 26.885 83.545 27.145 ;
        RECT 83.645 26.885 83.905 27.145 ;
        RECT 84.005 26.885 84.265 27.145 ;
        RECT 84.365 26.885 84.625 27.145 ;
        RECT 84.725 26.885 84.985 27.145 ;
        RECT 85.085 26.885 85.345 27.145 ;
        RECT 85.445 26.885 85.705 27.145 ;
        RECT 85.805 26.885 86.065 27.145 ;
        RECT 86.165 26.885 86.425 27.145 ;
        RECT 86.525 26.885 86.785 27.145 ;
        RECT 86.885 26.885 87.145 27.145 ;
        RECT 87.245 26.885 87.505 27.145 ;
        RECT 87.605 26.885 87.865 27.145 ;
        RECT 87.965 26.885 88.225 27.145 ;
        RECT 88.325 26.885 88.585 27.145 ;
        RECT 88.685 26.885 88.945 27.145 ;
        RECT 89.045 26.885 89.305 27.145 ;
        RECT 89.405 26.885 89.665 27.145 ;
        RECT 89.765 26.885 90.025 27.145 ;
        RECT 90.125 26.885 90.385 27.145 ;
        RECT 90.485 26.885 90.745 27.145 ;
        RECT 90.845 26.885 91.105 27.145 ;
        RECT 91.205 26.885 91.465 27.145 ;
        RECT 91.565 26.885 91.825 27.145 ;
        RECT 91.925 26.885 92.185 27.145 ;
        RECT 92.285 26.885 92.545 27.145 ;
        RECT 92.645 26.885 92.905 27.145 ;
        RECT 93.005 26.885 93.265 27.145 ;
        RECT 93.365 26.885 93.625 27.145 ;
        RECT 93.725 26.885 93.985 27.145 ;
        RECT 94.085 26.885 94.345 27.145 ;
        RECT 94.445 26.885 94.705 27.145 ;
        RECT 94.805 26.885 95.065 27.145 ;
        RECT 95.165 26.885 95.425 27.145 ;
        RECT 95.525 26.885 95.785 27.145 ;
        RECT 95.885 26.885 96.145 27.145 ;
        RECT 96.245 26.885 96.505 27.145 ;
        RECT 96.605 26.885 96.865 27.145 ;
        RECT 96.965 26.885 97.225 27.145 ;
        RECT 97.325 26.885 97.585 27.145 ;
        RECT 97.685 26.885 97.945 27.145 ;
        RECT 98.045 26.885 98.305 27.145 ;
        RECT 98.405 26.885 98.665 27.145 ;
        RECT 98.765 26.885 99.025 27.145 ;
        RECT 99.125 26.885 99.385 27.145 ;
        RECT 99.485 26.885 99.745 27.145 ;
        RECT 99.845 26.885 100.105 27.145 ;
        RECT 100.205 26.885 100.465 27.145 ;
        RECT 100.565 26.885 100.825 27.145 ;
        RECT 100.925 26.885 101.185 27.145 ;
        RECT 101.285 26.885 101.545 27.145 ;
        RECT 101.645 26.885 101.905 27.145 ;
        RECT 102.005 26.885 102.265 27.145 ;
        RECT 102.365 26.885 102.625 27.145 ;
        RECT 102.725 26.885 102.985 27.145 ;
        RECT 103.085 26.885 103.345 27.145 ;
        RECT 103.445 26.885 103.705 27.145 ;
        RECT 103.805 26.885 104.065 27.145 ;
        RECT 104.165 26.885 104.425 27.145 ;
        RECT 104.525 26.885 104.785 27.145 ;
        RECT 104.885 26.885 105.145 27.145 ;
        RECT 105.245 26.885 105.505 27.145 ;
        RECT 105.605 26.885 105.865 27.145 ;
        RECT 105.965 26.885 106.225 27.145 ;
        RECT 22.580 25.170 22.840 25.430 ;
        RECT 22.940 25.170 23.200 25.430 ;
        RECT 23.300 25.170 23.560 25.430 ;
        RECT 22.580 24.810 22.840 25.070 ;
        RECT 22.940 24.810 23.200 25.070 ;
        RECT 23.300 24.810 23.560 25.070 ;
        RECT 22.580 24.450 22.840 24.710 ;
        RECT 22.940 24.450 23.200 24.710 ;
        RECT 23.300 24.450 23.560 24.710 ;
        RECT 22.580 24.090 22.840 24.350 ;
        RECT 22.940 24.090 23.200 24.350 ;
        RECT 23.300 24.090 23.560 24.350 ;
        RECT 22.580 23.730 22.840 23.990 ;
        RECT 22.940 23.730 23.200 23.990 ;
        RECT 23.300 23.730 23.560 23.990 ;
        RECT 22.580 23.370 22.840 23.630 ;
        RECT 22.940 23.370 23.200 23.630 ;
        RECT 23.300 23.370 23.560 23.630 ;
        RECT 22.580 23.010 22.840 23.270 ;
        RECT 22.940 23.010 23.200 23.270 ;
        RECT 23.300 23.010 23.560 23.270 ;
        RECT 22.580 22.650 22.840 22.910 ;
        RECT 22.940 22.650 23.200 22.910 ;
        RECT 23.300 22.650 23.560 22.910 ;
        RECT 22.580 22.290 22.840 22.550 ;
        RECT 22.940 22.290 23.200 22.550 ;
        RECT 23.300 22.290 23.560 22.550 ;
        RECT 22.580 21.930 22.840 22.190 ;
        RECT 22.940 21.930 23.200 22.190 ;
        RECT 23.300 21.930 23.560 22.190 ;
        RECT 22.580 21.570 22.840 21.830 ;
        RECT 22.940 21.570 23.200 21.830 ;
        RECT 23.300 21.570 23.560 21.830 ;
        RECT 22.580 21.210 22.840 21.470 ;
        RECT 22.940 21.210 23.200 21.470 ;
        RECT 23.300 21.210 23.560 21.470 ;
        RECT 22.580 20.850 22.840 21.110 ;
        RECT 22.940 20.850 23.200 21.110 ;
        RECT 23.300 20.850 23.560 21.110 ;
        RECT 22.580 20.490 22.840 20.750 ;
        RECT 22.940 20.490 23.200 20.750 ;
        RECT 23.300 20.490 23.560 20.750 ;
        RECT 22.580 20.130 22.840 20.390 ;
        RECT 22.940 20.130 23.200 20.390 ;
        RECT 23.300 20.130 23.560 20.390 ;
        RECT 22.580 19.770 22.840 20.030 ;
        RECT 22.940 19.770 23.200 20.030 ;
        RECT 23.300 19.770 23.560 20.030 ;
        RECT 22.580 19.410 22.840 19.670 ;
        RECT 22.940 19.410 23.200 19.670 ;
        RECT 23.300 19.410 23.560 19.670 ;
        RECT 22.580 19.050 22.840 19.310 ;
        RECT 22.940 19.050 23.200 19.310 ;
        RECT 23.300 19.050 23.560 19.310 ;
        RECT 22.580 18.690 22.840 18.950 ;
        RECT 22.940 18.690 23.200 18.950 ;
        RECT 23.300 18.690 23.560 18.950 ;
        RECT 22.580 18.330 22.840 18.590 ;
        RECT 22.940 18.330 23.200 18.590 ;
        RECT 23.300 18.330 23.560 18.590 ;
        RECT 22.580 17.970 22.840 18.230 ;
        RECT 22.940 17.970 23.200 18.230 ;
        RECT 23.300 17.970 23.560 18.230 ;
        RECT 22.580 17.610 22.840 17.870 ;
        RECT 22.940 17.610 23.200 17.870 ;
        RECT 23.300 17.610 23.560 17.870 ;
        RECT 22.580 17.250 22.840 17.510 ;
        RECT 22.940 17.250 23.200 17.510 ;
        RECT 23.300 17.250 23.560 17.510 ;
        RECT 26.150 18.010 26.410 18.270 ;
        RECT 26.510 18.010 26.770 18.270 ;
        RECT 26.870 18.010 27.130 18.270 ;
        RECT 27.230 18.010 27.490 18.270 ;
        RECT 27.590 18.010 27.850 18.270 ;
        RECT 27.950 18.010 28.210 18.270 ;
        RECT 28.310 18.010 28.570 18.270 ;
        RECT 28.670 18.010 28.930 18.270 ;
        RECT 29.030 18.010 29.290 18.270 ;
        RECT 29.390 18.010 29.650 18.270 ;
        RECT 29.750 18.010 30.010 18.270 ;
        RECT 30.110 18.010 30.370 18.270 ;
        RECT 30.470 18.010 30.730 18.270 ;
        RECT 30.830 18.010 31.090 18.270 ;
        RECT 31.190 18.010 31.450 18.270 ;
        RECT 31.550 18.010 31.810 18.270 ;
        RECT 31.910 18.010 32.170 18.270 ;
        RECT 32.270 18.010 32.530 18.270 ;
        RECT 32.630 18.010 32.890 18.270 ;
        RECT 32.990 18.010 33.250 18.270 ;
        RECT 33.350 18.010 33.610 18.270 ;
        RECT 33.710 18.010 33.970 18.270 ;
        RECT 34.070 18.010 34.330 18.270 ;
        RECT 34.430 18.010 34.690 18.270 ;
        RECT 34.790 18.010 35.050 18.270 ;
        RECT 35.150 18.010 35.410 18.270 ;
        RECT 35.510 18.010 35.770 18.270 ;
        RECT 35.870 18.010 36.130 18.270 ;
        RECT 36.230 18.010 36.490 18.270 ;
        RECT 36.590 18.010 36.850 18.270 ;
        RECT 36.950 18.010 37.210 18.270 ;
        RECT 37.310 18.010 37.570 18.270 ;
        RECT 37.670 18.010 37.930 18.270 ;
        RECT 38.030 18.010 38.290 18.270 ;
        RECT 38.390 18.010 38.650 18.270 ;
        RECT 38.750 18.010 39.010 18.270 ;
        RECT 39.110 18.010 39.370 18.270 ;
        RECT 39.470 18.010 39.730 18.270 ;
        RECT 39.830 18.010 40.090 18.270 ;
        RECT 40.190 18.010 40.450 18.270 ;
        RECT 40.550 18.010 40.810 18.270 ;
        RECT 40.910 18.010 41.170 18.270 ;
        RECT 41.270 18.010 41.530 18.270 ;
        RECT 41.630 18.010 41.890 18.270 ;
        RECT 41.990 18.010 42.250 18.270 ;
        RECT 42.350 18.010 42.610 18.270 ;
        RECT 42.710 18.010 42.970 18.270 ;
        RECT 43.070 18.010 43.330 18.270 ;
        RECT 43.430 18.010 43.690 18.270 ;
        RECT 43.790 18.010 44.050 18.270 ;
        RECT 44.150 18.010 44.410 18.270 ;
        RECT 44.510 18.010 44.770 18.270 ;
        RECT 44.870 18.010 45.130 18.270 ;
        RECT 45.230 18.010 45.490 18.270 ;
        RECT 45.590 18.010 45.850 18.270 ;
        RECT 45.950 18.010 46.210 18.270 ;
        RECT 46.310 18.010 46.570 18.270 ;
        RECT 46.670 18.010 46.930 18.270 ;
        RECT 47.030 18.010 47.290 18.270 ;
        RECT 47.390 18.010 47.650 18.270 ;
        RECT 47.750 18.010 48.010 18.270 ;
        RECT 48.110 18.010 48.370 18.270 ;
        RECT 48.470 18.010 48.730 18.270 ;
        RECT 48.830 18.010 49.090 18.270 ;
        RECT 49.190 18.010 49.450 18.270 ;
        RECT 49.550 18.010 49.810 18.270 ;
        RECT 49.910 18.010 50.170 18.270 ;
        RECT 50.270 18.010 50.530 18.270 ;
        RECT 50.630 18.010 50.890 18.270 ;
        RECT 50.990 18.010 51.250 18.270 ;
        RECT 51.350 18.010 51.610 18.270 ;
        RECT 51.710 18.010 51.970 18.270 ;
        RECT 52.070 18.010 52.330 18.270 ;
        RECT 52.430 18.010 52.690 18.270 ;
        RECT 52.790 18.010 53.050 18.270 ;
        RECT 53.150 18.010 53.410 18.270 ;
        RECT 53.510 18.010 53.770 18.270 ;
        RECT 53.870 18.010 54.130 18.270 ;
        RECT 54.230 18.010 54.490 18.270 ;
        RECT 54.590 18.010 54.850 18.270 ;
        RECT 54.950 18.010 55.210 18.270 ;
        RECT 55.310 18.010 55.570 18.270 ;
        RECT 55.670 18.010 55.930 18.270 ;
        RECT 56.030 18.010 56.290 18.270 ;
        RECT 56.390 18.010 56.650 18.270 ;
        RECT 56.750 18.010 57.010 18.270 ;
        RECT 57.110 18.010 57.370 18.270 ;
        RECT 57.470 18.010 57.730 18.270 ;
        RECT 57.830 18.010 58.090 18.270 ;
        RECT 58.190 18.010 58.450 18.270 ;
        RECT 58.550 18.010 58.810 18.270 ;
        RECT 58.910 18.010 59.170 18.270 ;
        RECT 59.270 18.010 59.530 18.270 ;
        RECT 59.630 18.010 59.890 18.270 ;
        RECT 59.990 18.010 60.250 18.270 ;
        RECT 60.350 18.010 60.610 18.270 ;
        RECT 60.710 18.010 60.970 18.270 ;
        RECT 61.070 18.010 61.330 18.270 ;
        RECT 61.430 18.010 61.690 18.270 ;
        RECT 61.790 18.010 62.050 18.270 ;
        RECT 62.150 18.010 62.410 18.270 ;
        RECT 62.510 18.010 62.770 18.270 ;
        RECT 62.870 18.010 63.130 18.270 ;
        RECT 63.230 18.010 63.490 18.270 ;
        RECT 63.590 18.010 63.850 18.270 ;
        RECT 63.950 18.010 64.210 18.270 ;
        RECT 64.310 18.010 64.570 18.270 ;
        RECT 64.670 18.010 64.930 18.270 ;
        RECT 65.030 18.010 65.290 18.270 ;
        RECT 65.390 18.010 65.650 18.270 ;
        RECT 65.750 18.010 66.010 18.270 ;
        RECT 26.150 17.650 26.410 17.910 ;
        RECT 26.510 17.650 26.770 17.910 ;
        RECT 26.870 17.650 27.130 17.910 ;
        RECT 27.230 17.650 27.490 17.910 ;
        RECT 27.590 17.650 27.850 17.910 ;
        RECT 27.950 17.650 28.210 17.910 ;
        RECT 28.310 17.650 28.570 17.910 ;
        RECT 28.670 17.650 28.930 17.910 ;
        RECT 29.030 17.650 29.290 17.910 ;
        RECT 29.390 17.650 29.650 17.910 ;
        RECT 29.750 17.650 30.010 17.910 ;
        RECT 30.110 17.650 30.370 17.910 ;
        RECT 30.470 17.650 30.730 17.910 ;
        RECT 30.830 17.650 31.090 17.910 ;
        RECT 31.190 17.650 31.450 17.910 ;
        RECT 31.550 17.650 31.810 17.910 ;
        RECT 31.910 17.650 32.170 17.910 ;
        RECT 32.270 17.650 32.530 17.910 ;
        RECT 32.630 17.650 32.890 17.910 ;
        RECT 32.990 17.650 33.250 17.910 ;
        RECT 33.350 17.650 33.610 17.910 ;
        RECT 33.710 17.650 33.970 17.910 ;
        RECT 34.070 17.650 34.330 17.910 ;
        RECT 34.430 17.650 34.690 17.910 ;
        RECT 34.790 17.650 35.050 17.910 ;
        RECT 35.150 17.650 35.410 17.910 ;
        RECT 35.510 17.650 35.770 17.910 ;
        RECT 35.870 17.650 36.130 17.910 ;
        RECT 36.230 17.650 36.490 17.910 ;
        RECT 36.590 17.650 36.850 17.910 ;
        RECT 36.950 17.650 37.210 17.910 ;
        RECT 37.310 17.650 37.570 17.910 ;
        RECT 37.670 17.650 37.930 17.910 ;
        RECT 38.030 17.650 38.290 17.910 ;
        RECT 38.390 17.650 38.650 17.910 ;
        RECT 38.750 17.650 39.010 17.910 ;
        RECT 39.110 17.650 39.370 17.910 ;
        RECT 39.470 17.650 39.730 17.910 ;
        RECT 39.830 17.650 40.090 17.910 ;
        RECT 40.190 17.650 40.450 17.910 ;
        RECT 40.550 17.650 40.810 17.910 ;
        RECT 40.910 17.650 41.170 17.910 ;
        RECT 41.270 17.650 41.530 17.910 ;
        RECT 41.630 17.650 41.890 17.910 ;
        RECT 41.990 17.650 42.250 17.910 ;
        RECT 42.350 17.650 42.610 17.910 ;
        RECT 42.710 17.650 42.970 17.910 ;
        RECT 43.070 17.650 43.330 17.910 ;
        RECT 43.430 17.650 43.690 17.910 ;
        RECT 43.790 17.650 44.050 17.910 ;
        RECT 44.150 17.650 44.410 17.910 ;
        RECT 44.510 17.650 44.770 17.910 ;
        RECT 44.870 17.650 45.130 17.910 ;
        RECT 45.230 17.650 45.490 17.910 ;
        RECT 45.590 17.650 45.850 17.910 ;
        RECT 45.950 17.650 46.210 17.910 ;
        RECT 46.310 17.650 46.570 17.910 ;
        RECT 46.670 17.650 46.930 17.910 ;
        RECT 47.030 17.650 47.290 17.910 ;
        RECT 47.390 17.650 47.650 17.910 ;
        RECT 47.750 17.650 48.010 17.910 ;
        RECT 48.110 17.650 48.370 17.910 ;
        RECT 48.470 17.650 48.730 17.910 ;
        RECT 48.830 17.650 49.090 17.910 ;
        RECT 49.190 17.650 49.450 17.910 ;
        RECT 49.550 17.650 49.810 17.910 ;
        RECT 49.910 17.650 50.170 17.910 ;
        RECT 50.270 17.650 50.530 17.910 ;
        RECT 50.630 17.650 50.890 17.910 ;
        RECT 50.990 17.650 51.250 17.910 ;
        RECT 51.350 17.650 51.610 17.910 ;
        RECT 51.710 17.650 51.970 17.910 ;
        RECT 52.070 17.650 52.330 17.910 ;
        RECT 52.430 17.650 52.690 17.910 ;
        RECT 52.790 17.650 53.050 17.910 ;
        RECT 53.150 17.650 53.410 17.910 ;
        RECT 53.510 17.650 53.770 17.910 ;
        RECT 53.870 17.650 54.130 17.910 ;
        RECT 54.230 17.650 54.490 17.910 ;
        RECT 54.590 17.650 54.850 17.910 ;
        RECT 54.950 17.650 55.210 17.910 ;
        RECT 55.310 17.650 55.570 17.910 ;
        RECT 55.670 17.650 55.930 17.910 ;
        RECT 56.030 17.650 56.290 17.910 ;
        RECT 56.390 17.650 56.650 17.910 ;
        RECT 56.750 17.650 57.010 17.910 ;
        RECT 57.110 17.650 57.370 17.910 ;
        RECT 57.470 17.650 57.730 17.910 ;
        RECT 57.830 17.650 58.090 17.910 ;
        RECT 58.190 17.650 58.450 17.910 ;
        RECT 58.550 17.650 58.810 17.910 ;
        RECT 58.910 17.650 59.170 17.910 ;
        RECT 59.270 17.650 59.530 17.910 ;
        RECT 59.630 17.650 59.890 17.910 ;
        RECT 59.990 17.650 60.250 17.910 ;
        RECT 60.350 17.650 60.610 17.910 ;
        RECT 60.710 17.650 60.970 17.910 ;
        RECT 61.070 17.650 61.330 17.910 ;
        RECT 61.430 17.650 61.690 17.910 ;
        RECT 61.790 17.650 62.050 17.910 ;
        RECT 62.150 17.650 62.410 17.910 ;
        RECT 62.510 17.650 62.770 17.910 ;
        RECT 62.870 17.650 63.130 17.910 ;
        RECT 63.230 17.650 63.490 17.910 ;
        RECT 63.590 17.650 63.850 17.910 ;
        RECT 63.950 17.650 64.210 17.910 ;
        RECT 64.310 17.650 64.570 17.910 ;
        RECT 64.670 17.650 64.930 17.910 ;
        RECT 65.030 17.650 65.290 17.910 ;
        RECT 65.390 17.650 65.650 17.910 ;
        RECT 65.750 17.650 66.010 17.910 ;
        RECT 22.580 16.890 22.840 17.150 ;
        RECT 22.940 16.890 23.200 17.150 ;
        RECT 23.300 16.890 23.560 17.150 ;
        RECT 22.580 16.530 22.840 16.790 ;
        RECT 22.940 16.530 23.200 16.790 ;
        RECT 23.300 16.530 23.560 16.790 ;
        RECT 22.580 16.170 22.840 16.430 ;
        RECT 22.940 16.170 23.200 16.430 ;
        RECT 23.300 16.170 23.560 16.430 ;
        RECT 26.150 17.290 26.410 17.550 ;
        RECT 26.510 17.290 26.770 17.550 ;
        RECT 26.870 17.290 27.130 17.550 ;
        RECT 27.230 17.290 27.490 17.550 ;
        RECT 27.590 17.290 27.850 17.550 ;
        RECT 27.950 17.290 28.210 17.550 ;
        RECT 28.310 17.290 28.570 17.550 ;
        RECT 28.670 17.290 28.930 17.550 ;
        RECT 29.030 17.290 29.290 17.550 ;
        RECT 29.390 17.290 29.650 17.550 ;
        RECT 29.750 17.290 30.010 17.550 ;
        RECT 30.110 17.290 30.370 17.550 ;
        RECT 30.470 17.290 30.730 17.550 ;
        RECT 30.830 17.290 31.090 17.550 ;
        RECT 31.190 17.290 31.450 17.550 ;
        RECT 31.550 17.290 31.810 17.550 ;
        RECT 31.910 17.290 32.170 17.550 ;
        RECT 32.270 17.290 32.530 17.550 ;
        RECT 32.630 17.290 32.890 17.550 ;
        RECT 32.990 17.290 33.250 17.550 ;
        RECT 33.350 17.290 33.610 17.550 ;
        RECT 33.710 17.290 33.970 17.550 ;
        RECT 34.070 17.290 34.330 17.550 ;
        RECT 34.430 17.290 34.690 17.550 ;
        RECT 34.790 17.290 35.050 17.550 ;
        RECT 35.150 17.290 35.410 17.550 ;
        RECT 35.510 17.290 35.770 17.550 ;
        RECT 35.870 17.290 36.130 17.550 ;
        RECT 36.230 17.290 36.490 17.550 ;
        RECT 36.590 17.290 36.850 17.550 ;
        RECT 36.950 17.290 37.210 17.550 ;
        RECT 37.310 17.290 37.570 17.550 ;
        RECT 37.670 17.290 37.930 17.550 ;
        RECT 38.030 17.290 38.290 17.550 ;
        RECT 38.390 17.290 38.650 17.550 ;
        RECT 38.750 17.290 39.010 17.550 ;
        RECT 39.110 17.290 39.370 17.550 ;
        RECT 39.470 17.290 39.730 17.550 ;
        RECT 39.830 17.290 40.090 17.550 ;
        RECT 40.190 17.290 40.450 17.550 ;
        RECT 40.550 17.290 40.810 17.550 ;
        RECT 40.910 17.290 41.170 17.550 ;
        RECT 41.270 17.290 41.530 17.550 ;
        RECT 41.630 17.290 41.890 17.550 ;
        RECT 41.990 17.290 42.250 17.550 ;
        RECT 42.350 17.290 42.610 17.550 ;
        RECT 42.710 17.290 42.970 17.550 ;
        RECT 43.070 17.290 43.330 17.550 ;
        RECT 43.430 17.290 43.690 17.550 ;
        RECT 43.790 17.290 44.050 17.550 ;
        RECT 44.150 17.290 44.410 17.550 ;
        RECT 44.510 17.290 44.770 17.550 ;
        RECT 44.870 17.290 45.130 17.550 ;
        RECT 45.230 17.290 45.490 17.550 ;
        RECT 45.590 17.290 45.850 17.550 ;
        RECT 45.950 17.290 46.210 17.550 ;
        RECT 46.310 17.290 46.570 17.550 ;
        RECT 46.670 17.290 46.930 17.550 ;
        RECT 47.030 17.290 47.290 17.550 ;
        RECT 47.390 17.290 47.650 17.550 ;
        RECT 47.750 17.290 48.010 17.550 ;
        RECT 48.110 17.290 48.370 17.550 ;
        RECT 48.470 17.290 48.730 17.550 ;
        RECT 48.830 17.290 49.090 17.550 ;
        RECT 49.190 17.290 49.450 17.550 ;
        RECT 49.550 17.290 49.810 17.550 ;
        RECT 49.910 17.290 50.170 17.550 ;
        RECT 50.270 17.290 50.530 17.550 ;
        RECT 50.630 17.290 50.890 17.550 ;
        RECT 50.990 17.290 51.250 17.550 ;
        RECT 51.350 17.290 51.610 17.550 ;
        RECT 51.710 17.290 51.970 17.550 ;
        RECT 52.070 17.290 52.330 17.550 ;
        RECT 52.430 17.290 52.690 17.550 ;
        RECT 52.790 17.290 53.050 17.550 ;
        RECT 53.150 17.290 53.410 17.550 ;
        RECT 53.510 17.290 53.770 17.550 ;
        RECT 53.870 17.290 54.130 17.550 ;
        RECT 54.230 17.290 54.490 17.550 ;
        RECT 54.590 17.290 54.850 17.550 ;
        RECT 54.950 17.290 55.210 17.550 ;
        RECT 55.310 17.290 55.570 17.550 ;
        RECT 55.670 17.290 55.930 17.550 ;
        RECT 56.030 17.290 56.290 17.550 ;
        RECT 56.390 17.290 56.650 17.550 ;
        RECT 56.750 17.290 57.010 17.550 ;
        RECT 57.110 17.290 57.370 17.550 ;
        RECT 57.470 17.290 57.730 17.550 ;
        RECT 57.830 17.290 58.090 17.550 ;
        RECT 58.190 17.290 58.450 17.550 ;
        RECT 58.550 17.290 58.810 17.550 ;
        RECT 58.910 17.290 59.170 17.550 ;
        RECT 59.270 17.290 59.530 17.550 ;
        RECT 59.630 17.290 59.890 17.550 ;
        RECT 59.990 17.290 60.250 17.550 ;
        RECT 60.350 17.290 60.610 17.550 ;
        RECT 60.710 17.290 60.970 17.550 ;
        RECT 61.070 17.290 61.330 17.550 ;
        RECT 61.430 17.290 61.690 17.550 ;
        RECT 61.790 17.290 62.050 17.550 ;
        RECT 62.150 17.290 62.410 17.550 ;
        RECT 62.510 17.290 62.770 17.550 ;
        RECT 62.870 17.290 63.130 17.550 ;
        RECT 63.230 17.290 63.490 17.550 ;
        RECT 63.590 17.290 63.850 17.550 ;
        RECT 63.950 17.290 64.210 17.550 ;
        RECT 64.310 17.290 64.570 17.550 ;
        RECT 64.670 17.290 64.930 17.550 ;
        RECT 65.030 17.290 65.290 17.550 ;
        RECT 65.390 17.290 65.650 17.550 ;
        RECT 65.750 17.290 66.010 17.550 ;
        RECT 22.580 15.810 22.840 16.070 ;
        RECT 22.940 15.810 23.200 16.070 ;
        RECT 23.300 15.810 23.560 16.070 ;
        RECT 22.580 15.450 22.840 15.710 ;
        RECT 22.940 15.450 23.200 15.710 ;
        RECT 23.300 15.450 23.560 15.710 ;
        RECT 22.580 15.090 22.840 15.350 ;
        RECT 22.940 15.090 23.200 15.350 ;
        RECT 23.300 15.090 23.560 15.350 ;
        RECT 22.580 14.730 22.840 14.990 ;
        RECT 22.940 14.730 23.200 14.990 ;
        RECT 23.300 14.730 23.560 14.990 ;
        RECT 22.580 14.370 22.840 14.630 ;
        RECT 22.940 14.370 23.200 14.630 ;
        RECT 23.300 14.370 23.560 14.630 ;
        RECT 22.580 14.010 22.840 14.270 ;
        RECT 22.940 14.010 23.200 14.270 ;
        RECT 23.300 14.010 23.560 14.270 ;
        RECT 22.580 13.650 22.840 13.910 ;
        RECT 22.940 13.650 23.200 13.910 ;
        RECT 23.300 13.650 23.560 13.910 ;
        RECT 22.580 13.290 22.840 13.550 ;
        RECT 22.940 13.290 23.200 13.550 ;
        RECT 23.300 13.290 23.560 13.550 ;
        RECT 22.580 12.930 22.840 13.190 ;
        RECT 22.940 12.930 23.200 13.190 ;
        RECT 23.300 12.930 23.560 13.190 ;
        RECT 22.580 12.570 22.840 12.830 ;
        RECT 22.940 12.570 23.200 12.830 ;
        RECT 23.300 12.570 23.560 12.830 ;
        RECT 22.580 12.210 22.840 12.470 ;
        RECT 22.940 12.210 23.200 12.470 ;
        RECT 23.300 12.210 23.560 12.470 ;
        RECT 22.580 11.850 22.840 12.110 ;
        RECT 22.940 11.850 23.200 12.110 ;
        RECT 23.300 11.850 23.560 12.110 ;
        RECT 22.580 11.490 22.840 11.750 ;
        RECT 22.940 11.490 23.200 11.750 ;
        RECT 23.300 11.490 23.560 11.750 ;
        RECT 22.580 11.130 22.840 11.390 ;
        RECT 22.940 11.130 23.200 11.390 ;
        RECT 23.300 11.130 23.560 11.390 ;
        RECT 22.580 10.770 22.840 11.030 ;
        RECT 22.940 10.770 23.200 11.030 ;
        RECT 23.300 10.770 23.560 11.030 ;
        RECT 22.580 10.410 22.840 10.670 ;
        RECT 22.940 10.410 23.200 10.670 ;
        RECT 23.300 10.410 23.560 10.670 ;
        RECT 22.580 10.050 22.840 10.310 ;
        RECT 22.940 10.050 23.200 10.310 ;
        RECT 23.300 10.050 23.560 10.310 ;
        RECT 22.580 9.690 22.840 9.950 ;
        RECT 22.940 9.690 23.200 9.950 ;
        RECT 23.300 9.690 23.560 9.950 ;
        RECT 22.580 9.330 22.840 9.590 ;
        RECT 22.940 9.330 23.200 9.590 ;
        RECT 23.300 9.330 23.560 9.590 ;
        RECT 22.580 8.970 22.840 9.230 ;
        RECT 22.940 8.970 23.200 9.230 ;
        RECT 23.300 8.970 23.560 9.230 ;
        RECT 22.580 8.610 22.840 8.870 ;
        RECT 22.940 8.610 23.200 8.870 ;
        RECT 23.300 8.610 23.560 8.870 ;
        RECT 22.580 8.250 22.840 8.510 ;
        RECT 22.940 8.250 23.200 8.510 ;
        RECT 23.300 8.250 23.560 8.510 ;
        RECT 22.580 7.890 22.840 8.150 ;
        RECT 22.940 7.890 23.200 8.150 ;
        RECT 23.300 7.890 23.560 8.150 ;
        RECT 22.580 7.530 22.840 7.790 ;
        RECT 22.940 7.530 23.200 7.790 ;
        RECT 23.300 7.530 23.560 7.790 ;
        RECT 22.580 7.170 22.840 7.430 ;
        RECT 22.940 7.170 23.200 7.430 ;
        RECT 23.300 7.170 23.560 7.430 ;
        RECT 22.580 6.810 22.840 7.070 ;
        RECT 22.940 6.810 23.200 7.070 ;
        RECT 23.300 6.810 23.560 7.070 ;
        RECT 22.580 6.450 22.840 6.710 ;
        RECT 22.940 6.450 23.200 6.710 ;
        RECT 23.300 6.450 23.560 6.710 ;
        RECT 22.580 6.090 22.840 6.350 ;
        RECT 22.940 6.090 23.200 6.350 ;
        RECT 23.300 6.090 23.560 6.350 ;
        RECT 22.580 5.730 22.840 5.990 ;
        RECT 22.940 5.730 23.200 5.990 ;
        RECT 23.300 5.730 23.560 5.990 ;
      LAYER met2 ;
        RECT 84.955 102.980 102.975 104.460 ;
        RECT 91.290 101.685 95.970 102.365 ;
        RECT 106.710 101.505 109.830 102.825 ;
        RECT 11.090 90.310 52.010 92.350 ;
        RECT 56.320 88.410 97.240 90.450 ;
        RECT 16.000 47.455 18.040 88.375 ;
        RECT 99.805 48.820 101.845 89.740 ;
        RECT 22.050 5.200 24.090 46.120 ;
        RECT 65.835 26.355 106.755 28.395 ;
        RECT 25.620 16.760 66.540 18.800 ;
      LAYER via2 ;
        RECT 85.630 103.580 85.910 103.860 ;
        RECT 86.030 103.580 86.310 103.860 ;
        RECT 86.430 103.580 86.710 103.860 ;
        RECT 86.830 103.580 87.110 103.860 ;
        RECT 87.230 103.580 87.510 103.860 ;
        RECT 87.630 103.580 87.910 103.860 ;
        RECT 88.030 103.580 88.310 103.860 ;
        RECT 88.430 103.580 88.710 103.860 ;
        RECT 88.830 103.580 89.110 103.860 ;
        RECT 89.230 103.580 89.510 103.860 ;
        RECT 89.630 103.580 89.910 103.860 ;
        RECT 90.030 103.580 90.310 103.860 ;
        RECT 90.430 103.580 90.710 103.860 ;
        RECT 90.830 103.580 91.110 103.860 ;
        RECT 91.230 103.580 91.510 103.860 ;
        RECT 91.630 103.580 91.910 103.860 ;
        RECT 92.030 103.580 92.310 103.860 ;
        RECT 92.430 103.580 92.710 103.860 ;
        RECT 92.830 103.580 93.110 103.860 ;
        RECT 93.230 103.580 93.510 103.860 ;
        RECT 93.630 103.580 93.910 103.860 ;
        RECT 94.030 103.580 94.310 103.860 ;
        RECT 94.430 103.580 94.710 103.860 ;
        RECT 94.830 103.580 95.110 103.860 ;
        RECT 95.230 103.580 95.510 103.860 ;
        RECT 95.630 103.580 95.910 103.860 ;
        RECT 96.030 103.580 96.310 103.860 ;
        RECT 96.430 103.580 96.710 103.860 ;
        RECT 96.830 103.580 97.110 103.860 ;
        RECT 97.230 103.580 97.510 103.860 ;
        RECT 97.630 103.580 97.910 103.860 ;
        RECT 98.030 103.580 98.310 103.860 ;
        RECT 98.430 103.580 98.710 103.860 ;
        RECT 98.830 103.580 99.110 103.860 ;
        RECT 99.230 103.580 99.510 103.860 ;
        RECT 99.630 103.580 99.910 103.860 ;
        RECT 100.030 103.580 100.310 103.860 ;
        RECT 100.430 103.580 100.710 103.860 ;
        RECT 100.830 103.580 101.110 103.860 ;
        RECT 101.230 103.580 101.510 103.860 ;
        RECT 101.630 103.580 101.910 103.860 ;
        RECT 102.030 103.580 102.310 103.860 ;
        RECT 107.230 102.025 107.510 102.305 ;
        RECT 107.680 102.025 107.960 102.305 ;
        RECT 108.130 102.025 108.410 102.305 ;
        RECT 108.580 102.025 108.860 102.305 ;
        RECT 109.030 102.025 109.310 102.305 ;
        RECT 11.830 90.990 51.310 91.670 ;
        RECT 57.040 89.090 96.520 89.770 ;
        RECT 16.680 48.175 17.360 87.655 ;
        RECT 100.485 49.540 101.165 89.020 ;
        RECT 22.730 5.920 23.410 45.400 ;
        RECT 66.555 27.035 106.035 27.715 ;
        RECT 26.340 17.440 65.820 18.120 ;
      LAYER met3 ;
        RECT 0.000 98.620 9.690 111.520 ;
        RECT 84.670 98.620 110.355 104.580 ;
        RECT 0.000 91.140 110.355 98.620 ;
        RECT 0.000 55.210 108.910 91.140 ;
        RECT 0.000 50.650 2.000 55.210 ;
        RECT 15.740 47.230 108.910 55.210 ;
        RECT 21.790 26.070 108.910 47.230 ;
        RECT 21.790 8.590 98.095 26.070 ;
        RECT 21.790 5.200 24.390 8.590 ;
        RECT 62.270 8.585 98.095 8.590 ;
      LAYER via3 ;
        RECT 0.240 51.000 1.760 111.320 ;
      LAYER met4 ;
        RECT 0.000 0.000 2.000 111.520 ;
    END
  END VPWR
  OBS
      LAYER pwell ;
        RECT 95.255 106.335 95.425 106.525 ;
        RECT 100.775 106.335 100.945 106.525 ;
        RECT 102.150 106.335 102.320 106.525 ;
        RECT 85.820 105.425 95.570 106.335 ;
        RECT 95.960 105.425 101.090 106.335 ;
        RECT 101.100 105.555 102.470 106.335 ;
        RECT 11.340 101.915 12.600 102.415 ;
        RECT 12.695 101.915 18.455 103.565 ;
      LAYER nwell ;
        RECT 85.265 103.530 102.665 105.135 ;
      LAYER pwell ;
        RECT 11.340 101.355 41.680 101.915 ;
        RECT 11.420 98.335 41.680 101.355 ;
        RECT 56.570 100.015 57.830 100.515 ;
        RECT 57.960 100.015 63.720 101.715 ;
        RECT 90.750 101.145 96.510 102.905 ;
        RECT 56.570 99.455 86.910 100.015 ;
        RECT 56.650 96.435 86.910 99.455 ;
        RECT 110.850 89.410 111.910 89.490 ;
        RECT 107.830 88.230 111.910 89.410 ;
        RECT 107.830 88.100 111.410 88.230 ;
        RECT 107.830 82.340 113.055 88.100 ;
        RECT 6.435 54.830 10.015 78.045 ;
        RECT 107.830 59.150 111.410 82.340 ;
        RECT 4.755 49.070 10.015 54.830 ;
        RECT 6.435 48.965 10.015 49.070 ;
        RECT 5.935 47.785 10.015 48.965 ;
        RECT 5.935 47.705 6.995 47.785 ;
        RECT 12.485 12.630 16.065 35.790 ;
        RECT 76.165 17.350 106.425 20.370 ;
        RECT 76.165 16.790 106.505 17.350 ;
        RECT 99.380 15.125 105.140 16.790 ;
        RECT 105.245 16.290 106.505 16.790 ;
        RECT 10.730 6.870 16.065 12.630 ;
        RECT 35.950 7.755 66.210 10.775 ;
        RECT 35.950 7.195 66.290 7.755 ;
        RECT 12.485 6.710 16.065 6.870 ;
        RECT 11.985 5.530 16.065 6.710 ;
        RECT 59.170 5.555 64.930 7.195 ;
        RECT 65.030 6.695 66.290 7.195 ;
        RECT 11.985 5.450 13.045 5.530 ;
      LAYER li1 ;
        RECT 117.035 107.070 119.215 107.420 ;
        RECT 119.615 107.070 121.795 107.420 ;
        RECT 93.050 105.705 93.380 106.180 ;
        RECT 93.890 105.705 94.220 106.180 ;
        RECT 94.730 105.705 95.060 106.180 ;
        RECT 92.710 105.535 95.060 105.705 ;
        RECT 96.550 105.705 96.720 106.185 ;
        RECT 97.390 105.705 97.560 106.185 ;
        RECT 98.230 105.705 98.400 106.185 ;
        RECT 99.070 105.705 99.240 106.185 ;
        RECT 99.910 105.705 100.080 106.180 ;
        RECT 100.750 105.705 100.920 106.185 ;
        RECT 96.550 105.535 99.240 105.705 ;
        RECT 99.500 105.535 100.920 105.705 ;
        RECT 101.180 105.680 101.440 106.185 ;
        RECT 102.130 105.805 102.300 106.185 ;
        RECT 92.710 105.365 92.885 105.535 ;
        RECT 96.550 105.365 96.805 105.535 ;
        RECT 99.500 105.365 99.675 105.535 ;
        RECT 101.180 105.365 101.360 105.680 ;
        RECT 101.635 105.635 102.300 105.805 ;
        RECT 114.550 105.800 116.730 106.150 ;
        RECT 122.100 105.800 124.280 106.150 ;
        RECT 101.635 105.380 101.805 105.635 ;
        RECT 86.165 105.165 92.885 105.365 ;
        RECT 93.090 105.165 96.805 105.365 ;
        RECT 97.050 105.195 99.675 105.365 ;
        RECT 92.710 104.995 92.885 105.165 ;
        RECT 96.550 104.995 96.805 105.165 ;
        RECT 99.500 104.995 99.675 105.195 ;
        RECT 99.855 105.165 101.360 105.365 ;
        RECT 92.710 104.825 95.060 104.995 ;
        RECT 93.050 103.975 93.380 104.825 ;
        RECT 93.890 103.975 94.220 104.825 ;
        RECT 94.730 103.975 95.060 104.825 ;
        RECT 96.550 104.825 99.240 104.995 ;
        RECT 99.500 104.825 101.000 104.995 ;
        RECT 96.550 103.975 96.720 104.825 ;
        RECT 97.390 103.975 97.560 104.825 ;
        RECT 98.230 103.975 98.400 104.825 ;
        RECT 99.070 103.975 99.240 104.825 ;
        RECT 99.830 103.975 100.160 104.825 ;
        RECT 100.670 103.975 101.000 104.825 ;
        RECT 101.180 104.880 101.360 105.165 ;
        RECT 101.530 105.050 101.805 105.380 ;
        RECT 102.030 105.085 102.690 105.455 ;
        RECT 101.635 104.905 101.805 105.050 ;
        RECT 139.585 105.005 140.475 105.595 ;
        RECT 101.180 103.975 101.450 104.880 ;
        RECT 101.635 104.735 102.310 104.905 ;
        RECT 102.130 103.975 102.310 104.735 ;
        RECT 112.065 104.530 114.245 104.880 ;
        RECT 124.585 104.530 126.765 104.880 ;
        RECT 109.580 103.260 111.760 103.610 ;
        RECT 127.070 103.260 129.250 103.610 ;
        RECT 13.275 102.785 13.475 102.985 ;
        RECT 13.675 102.785 13.875 102.985 ;
        RECT 14.075 102.785 14.275 102.985 ;
        RECT 14.475 102.785 14.675 102.985 ;
        RECT 14.875 102.785 15.075 102.985 ;
        RECT 15.275 102.785 15.475 102.985 ;
        RECT 15.675 102.785 15.875 102.985 ;
        RECT 16.075 102.785 16.275 102.985 ;
        RECT 16.475 102.785 16.675 102.985 ;
        RECT 16.875 102.785 17.075 102.985 ;
        RECT 17.275 102.785 17.475 102.985 ;
        RECT 17.675 102.785 17.875 102.985 ;
        RECT 13.275 102.385 13.475 102.585 ;
        RECT 13.675 102.385 13.875 102.585 ;
        RECT 14.075 102.385 14.275 102.585 ;
        RECT 14.475 102.385 14.675 102.585 ;
        RECT 14.875 102.385 15.075 102.585 ;
        RECT 15.275 102.385 15.475 102.585 ;
        RECT 15.675 102.385 15.875 102.585 ;
        RECT 16.075 102.385 16.275 102.585 ;
        RECT 16.475 102.385 16.675 102.585 ;
        RECT 16.875 102.385 17.075 102.585 ;
        RECT 17.275 102.385 17.475 102.585 ;
        RECT 17.675 102.385 17.875 102.585 ;
        RECT 136.390 102.450 136.560 102.620 ;
        RECT 91.330 102.125 91.530 102.325 ;
        RECT 91.730 102.125 91.930 102.325 ;
        RECT 92.130 102.125 92.330 102.325 ;
        RECT 92.530 102.125 92.730 102.325 ;
        RECT 92.930 102.125 93.130 102.325 ;
        RECT 93.330 102.125 93.530 102.325 ;
        RECT 93.730 102.125 93.930 102.325 ;
        RECT 94.130 102.125 94.330 102.325 ;
        RECT 94.530 102.125 94.730 102.325 ;
        RECT 94.930 102.125 95.130 102.325 ;
        RECT 95.330 102.125 95.530 102.325 ;
        RECT 95.730 102.125 95.930 102.325 ;
        RECT 11.020 101.720 11.190 102.050 ;
        RECT 109.580 101.990 111.760 102.340 ;
        RECT 112.160 101.990 114.340 102.340 ;
        RECT 114.550 101.990 116.730 102.340 ;
        RECT 117.130 101.990 119.310 102.340 ;
        RECT 119.520 101.990 121.700 102.340 ;
        RECT 122.100 101.990 124.280 102.340 ;
        RECT 124.490 101.990 126.670 102.340 ;
        RECT 127.070 101.990 129.250 102.340 ;
        RECT 91.330 101.725 91.530 101.925 ;
        RECT 91.730 101.725 91.930 101.925 ;
        RECT 92.130 101.725 92.330 101.925 ;
        RECT 92.530 101.725 92.730 101.925 ;
        RECT 92.930 101.725 93.130 101.925 ;
        RECT 93.330 101.725 93.530 101.925 ;
        RECT 93.730 101.725 93.930 101.925 ;
        RECT 94.130 101.725 94.330 101.925 ;
        RECT 94.530 101.725 94.730 101.925 ;
        RECT 94.930 101.725 95.130 101.925 ;
        RECT 95.330 101.725 95.530 101.925 ;
        RECT 95.730 101.725 95.930 101.925 ;
        RECT 11.625 101.190 41.475 101.720 ;
        RECT 11.100 99.240 11.270 101.010 ;
        RECT 58.540 100.935 58.740 101.135 ;
        RECT 58.940 100.935 59.140 101.135 ;
        RECT 59.340 100.935 59.540 101.135 ;
        RECT 59.740 100.935 59.940 101.135 ;
        RECT 60.140 100.935 60.340 101.135 ;
        RECT 60.540 100.935 60.740 101.135 ;
        RECT 60.940 100.935 61.140 101.135 ;
        RECT 61.340 100.935 61.540 101.135 ;
        RECT 61.740 100.935 61.940 101.135 ;
        RECT 62.140 100.935 62.340 101.135 ;
        RECT 62.540 100.935 62.740 101.135 ;
        RECT 62.940 100.935 63.140 101.135 ;
        RECT 58.540 100.535 58.740 100.735 ;
        RECT 58.940 100.535 59.140 100.735 ;
        RECT 59.340 100.535 59.540 100.735 ;
        RECT 59.740 100.535 59.940 100.735 ;
        RECT 60.140 100.535 60.340 100.735 ;
        RECT 60.540 100.535 60.740 100.735 ;
        RECT 60.940 100.535 61.140 100.735 ;
        RECT 61.340 100.535 61.540 100.735 ;
        RECT 61.740 100.535 61.940 100.735 ;
        RECT 62.140 100.535 62.340 100.735 ;
        RECT 62.540 100.535 62.740 100.735 ;
        RECT 62.940 100.535 63.140 100.735 ;
        RECT 109.675 100.720 111.855 101.070 ;
        RECT 112.065 100.720 114.245 101.070 ;
        RECT 114.645 100.720 116.825 101.070 ;
        RECT 117.035 100.720 119.215 101.070 ;
        RECT 119.615 100.720 121.795 101.070 ;
        RECT 122.005 100.720 124.185 101.070 ;
        RECT 124.585 100.720 126.765 101.070 ;
        RECT 126.975 100.720 129.155 101.070 ;
        RECT 56.250 99.820 56.420 100.150 ;
        RECT 56.855 99.290 86.705 99.820 ;
        RECT 11.625 98.530 41.475 99.060 ;
        RECT 11.585 97.080 51.515 97.970 ;
        RECT 56.330 97.340 56.500 99.110 ;
        RECT 11.100 93.050 11.270 96.980 ;
        RECT 56.855 96.630 86.705 97.160 ;
        RECT 56.815 95.180 96.745 96.070 ;
        RECT 56.330 91.150 56.500 95.080 ;
        RECT 102.545 89.560 106.475 89.730 ;
        RECT 108.735 89.560 110.505 89.730 ;
        RECT 111.215 89.640 111.545 89.810 ;
        RECT 5.335 54.050 5.535 54.250 ;
        RECT 5.735 54.050 5.935 54.250 ;
        RECT 5.335 53.650 5.535 53.850 ;
        RECT 5.735 53.650 5.935 53.850 ;
        RECT 5.335 53.250 5.535 53.450 ;
        RECT 5.735 53.250 5.935 53.450 ;
        RECT 5.335 52.850 5.535 53.050 ;
        RECT 5.735 52.850 5.935 53.050 ;
        RECT 5.335 52.450 5.535 52.650 ;
        RECT 5.735 52.450 5.935 52.650 ;
        RECT 5.335 52.050 5.535 52.250 ;
        RECT 5.735 52.050 5.935 52.250 ;
        RECT 5.335 51.650 5.535 51.850 ;
        RECT 5.735 51.650 5.935 51.850 ;
        RECT 5.335 51.250 5.535 51.450 ;
        RECT 5.735 51.250 5.935 51.450 ;
        RECT 5.335 50.850 5.535 51.050 ;
        RECT 5.735 50.850 5.935 51.050 ;
        RECT 5.335 50.450 5.535 50.650 ;
        RECT 5.735 50.450 5.935 50.650 ;
        RECT 5.335 50.050 5.535 50.250 ;
        RECT 5.735 50.050 5.935 50.250 ;
        RECT 5.335 49.650 5.535 49.850 ;
        RECT 5.735 49.650 5.935 49.850 ;
        RECT 6.630 47.990 7.160 77.840 ;
        RECT 9.290 47.990 9.820 77.840 ;
        RECT 10.380 47.950 11.270 87.880 ;
        RECT 106.575 49.315 107.465 89.245 ;
        RECT 108.025 59.355 108.555 89.205 ;
        RECT 110.685 59.355 111.215 89.205 ;
        RECT 111.875 87.320 112.075 87.520 ;
        RECT 112.275 87.320 112.475 87.520 ;
        RECT 111.875 86.920 112.075 87.120 ;
        RECT 112.275 86.920 112.475 87.120 ;
        RECT 111.875 86.520 112.075 86.720 ;
        RECT 112.275 86.520 112.475 86.720 ;
        RECT 111.875 86.120 112.075 86.320 ;
        RECT 112.275 86.120 112.475 86.320 ;
        RECT 111.875 85.720 112.075 85.920 ;
        RECT 112.275 85.720 112.475 85.920 ;
        RECT 111.875 85.320 112.075 85.520 ;
        RECT 112.275 85.320 112.475 85.520 ;
        RECT 111.875 84.920 112.075 85.120 ;
        RECT 112.275 84.920 112.475 85.120 ;
        RECT 111.875 84.520 112.075 84.720 ;
        RECT 112.275 84.520 112.475 84.720 ;
        RECT 111.875 84.120 112.075 84.320 ;
        RECT 112.275 84.120 112.475 84.320 ;
        RECT 111.875 83.720 112.075 83.920 ;
        RECT 112.275 83.720 112.475 83.920 ;
        RECT 111.875 83.320 112.075 83.520 ;
        RECT 112.275 83.320 112.475 83.520 ;
        RECT 111.875 82.920 112.075 83.120 ;
        RECT 112.275 82.920 112.475 83.120 ;
        RECT 6.300 47.385 6.630 47.555 ;
        RECT 7.340 47.465 9.110 47.635 ;
        RECT 11.370 47.465 15.300 47.635 ;
        RECT 11.310 11.850 11.510 12.050 ;
        RECT 11.710 11.850 11.910 12.050 ;
        RECT 11.310 11.450 11.510 11.650 ;
        RECT 11.710 11.450 11.910 11.650 ;
        RECT 11.310 11.050 11.510 11.250 ;
        RECT 11.710 11.050 11.910 11.250 ;
        RECT 11.310 10.650 11.510 10.850 ;
        RECT 11.710 10.650 11.910 10.850 ;
        RECT 11.310 10.250 11.510 10.450 ;
        RECT 11.710 10.250 11.910 10.450 ;
        RECT 11.310 9.850 11.510 10.050 ;
        RECT 11.710 9.850 11.910 10.050 ;
        RECT 11.310 9.450 11.510 9.650 ;
        RECT 11.710 9.450 11.910 9.650 ;
        RECT 11.310 9.050 11.510 9.250 ;
        RECT 11.710 9.050 11.910 9.250 ;
        RECT 11.310 8.650 11.510 8.850 ;
        RECT 11.710 8.650 11.910 8.850 ;
        RECT 11.310 8.250 11.510 8.450 ;
        RECT 11.710 8.250 11.910 8.450 ;
        RECT 11.310 7.850 11.510 8.050 ;
        RECT 11.710 7.850 11.910 8.050 ;
        RECT 11.310 7.450 11.510 7.650 ;
        RECT 11.710 7.450 11.910 7.650 ;
        RECT 12.680 5.735 13.210 35.585 ;
        RECT 15.340 5.735 15.870 35.585 ;
        RECT 16.430 5.695 17.320 45.625 ;
        RECT 106.575 21.725 106.745 25.655 ;
        RECT 66.330 20.735 106.260 21.625 ;
        RECT 76.370 19.645 106.220 20.175 ;
        RECT 106.575 17.695 106.745 19.465 ;
        RECT 76.370 16.985 106.220 17.515 ;
        RECT 106.655 16.655 106.825 16.985 ;
        RECT 99.960 16.105 100.160 16.305 ;
        RECT 100.360 16.105 100.560 16.305 ;
        RECT 100.760 16.105 100.960 16.305 ;
        RECT 101.160 16.105 101.360 16.305 ;
        RECT 101.560 16.105 101.760 16.305 ;
        RECT 101.960 16.105 102.160 16.305 ;
        RECT 102.360 16.105 102.560 16.305 ;
        RECT 102.760 16.105 102.960 16.305 ;
        RECT 103.160 16.105 103.360 16.305 ;
        RECT 103.560 16.105 103.760 16.305 ;
        RECT 103.960 16.105 104.160 16.305 ;
        RECT 104.360 16.105 104.560 16.305 ;
        RECT 66.360 12.130 66.530 16.060 ;
        RECT 99.960 15.705 100.160 15.905 ;
        RECT 100.360 15.705 100.560 15.905 ;
        RECT 100.760 15.705 100.960 15.905 ;
        RECT 101.160 15.705 101.360 15.905 ;
        RECT 101.560 15.705 101.760 15.905 ;
        RECT 101.960 15.705 102.160 15.905 ;
        RECT 102.360 15.705 102.560 15.905 ;
        RECT 102.760 15.705 102.960 15.905 ;
        RECT 103.160 15.705 103.360 15.905 ;
        RECT 103.560 15.705 103.760 15.905 ;
        RECT 103.960 15.705 104.160 15.905 ;
        RECT 104.360 15.705 104.560 15.905 ;
        RECT 26.115 11.140 66.045 12.030 ;
        RECT 36.155 10.050 66.005 10.580 ;
        RECT 66.360 8.100 66.530 9.870 ;
        RECT 36.155 7.390 66.005 7.920 ;
        RECT 66.440 7.060 66.610 7.390 ;
        RECT 59.750 6.535 59.950 6.735 ;
        RECT 60.150 6.535 60.350 6.735 ;
        RECT 60.550 6.535 60.750 6.735 ;
        RECT 60.950 6.535 61.150 6.735 ;
        RECT 61.350 6.535 61.550 6.735 ;
        RECT 61.750 6.535 61.950 6.735 ;
        RECT 62.150 6.535 62.350 6.735 ;
        RECT 62.550 6.535 62.750 6.735 ;
        RECT 62.950 6.535 63.150 6.735 ;
        RECT 63.350 6.535 63.550 6.735 ;
        RECT 63.750 6.535 63.950 6.735 ;
        RECT 64.150 6.535 64.350 6.735 ;
        RECT 59.750 6.135 59.950 6.335 ;
        RECT 60.150 6.135 60.350 6.335 ;
        RECT 60.550 6.135 60.750 6.335 ;
        RECT 60.950 6.135 61.150 6.335 ;
        RECT 61.350 6.135 61.550 6.335 ;
        RECT 61.750 6.135 61.950 6.335 ;
        RECT 62.150 6.135 62.350 6.335 ;
        RECT 62.550 6.135 62.750 6.335 ;
        RECT 62.950 6.135 63.150 6.335 ;
        RECT 63.350 6.135 63.550 6.335 ;
        RECT 63.750 6.135 63.950 6.335 ;
        RECT 64.150 6.135 64.350 6.335 ;
        RECT 12.350 5.130 12.680 5.300 ;
        RECT 13.390 5.210 15.160 5.380 ;
        RECT 17.420 5.210 21.350 5.380 ;
      LAYER mcon ;
        RECT 117.145 107.160 117.315 107.330 ;
        RECT 117.505 107.160 117.675 107.330 ;
        RECT 117.865 107.160 118.035 107.330 ;
        RECT 118.225 107.160 118.395 107.330 ;
        RECT 118.585 107.160 118.755 107.330 ;
        RECT 118.945 107.160 119.115 107.330 ;
        RECT 119.710 107.160 119.880 107.330 ;
        RECT 120.070 107.160 120.240 107.330 ;
        RECT 120.430 107.160 120.600 107.330 ;
        RECT 120.790 107.160 120.960 107.330 ;
        RECT 121.150 107.160 121.320 107.330 ;
        RECT 121.510 107.160 121.680 107.330 ;
        RECT 114.660 105.890 114.830 106.060 ;
        RECT 115.020 105.890 115.190 106.060 ;
        RECT 115.380 105.890 115.550 106.060 ;
        RECT 115.740 105.890 115.910 106.060 ;
        RECT 116.100 105.890 116.270 106.060 ;
        RECT 116.460 105.890 116.630 106.060 ;
        RECT 122.195 105.890 122.365 106.060 ;
        RECT 122.555 105.890 122.725 106.060 ;
        RECT 122.915 105.890 123.085 106.060 ;
        RECT 123.275 105.890 123.445 106.060 ;
        RECT 123.635 105.890 123.805 106.060 ;
        RECT 123.995 105.890 124.165 106.060 ;
        RECT 102.090 105.180 102.260 105.350 ;
        RECT 102.485 105.180 102.655 105.350 ;
        RECT 112.175 104.620 112.345 104.790 ;
        RECT 112.535 104.620 112.705 104.790 ;
        RECT 112.895 104.620 113.065 104.790 ;
        RECT 113.255 104.620 113.425 104.790 ;
        RECT 113.615 104.620 113.785 104.790 ;
        RECT 113.975 104.620 114.145 104.790 ;
        RECT 124.680 104.620 124.850 104.790 ;
        RECT 125.040 104.620 125.210 104.790 ;
        RECT 125.400 104.620 125.570 104.790 ;
        RECT 125.760 104.620 125.930 104.790 ;
        RECT 126.120 104.620 126.290 104.790 ;
        RECT 126.480 104.620 126.650 104.790 ;
        RECT 109.690 103.350 109.860 103.520 ;
        RECT 110.050 103.350 110.220 103.520 ;
        RECT 110.410 103.350 110.580 103.520 ;
        RECT 110.770 103.350 110.940 103.520 ;
        RECT 111.130 103.350 111.300 103.520 ;
        RECT 111.490 103.350 111.660 103.520 ;
        RECT 127.165 103.350 127.335 103.520 ;
        RECT 127.525 103.350 127.695 103.520 ;
        RECT 127.885 103.350 128.055 103.520 ;
        RECT 128.245 103.350 128.415 103.520 ;
        RECT 128.605 103.350 128.775 103.520 ;
        RECT 128.965 103.350 129.135 103.520 ;
        RECT 109.690 102.080 109.860 102.250 ;
        RECT 110.050 102.080 110.220 102.250 ;
        RECT 110.410 102.080 110.580 102.250 ;
        RECT 110.770 102.080 110.940 102.250 ;
        RECT 111.130 102.080 111.300 102.250 ;
        RECT 111.490 102.080 111.660 102.250 ;
        RECT 112.255 102.080 112.425 102.250 ;
        RECT 112.615 102.080 112.785 102.250 ;
        RECT 112.975 102.080 113.145 102.250 ;
        RECT 113.335 102.080 113.505 102.250 ;
        RECT 113.695 102.080 113.865 102.250 ;
        RECT 114.055 102.080 114.225 102.250 ;
        RECT 114.660 102.080 114.830 102.250 ;
        RECT 115.020 102.080 115.190 102.250 ;
        RECT 115.380 102.080 115.550 102.250 ;
        RECT 115.740 102.080 115.910 102.250 ;
        RECT 116.100 102.080 116.270 102.250 ;
        RECT 116.460 102.080 116.630 102.250 ;
        RECT 117.225 102.080 117.395 102.250 ;
        RECT 117.585 102.080 117.755 102.250 ;
        RECT 117.945 102.080 118.115 102.250 ;
        RECT 118.305 102.080 118.475 102.250 ;
        RECT 118.665 102.080 118.835 102.250 ;
        RECT 119.025 102.080 119.195 102.250 ;
        RECT 119.630 102.080 119.800 102.250 ;
        RECT 119.990 102.080 120.160 102.250 ;
        RECT 120.350 102.080 120.520 102.250 ;
        RECT 120.710 102.080 120.880 102.250 ;
        RECT 121.070 102.080 121.240 102.250 ;
        RECT 121.430 102.080 121.600 102.250 ;
        RECT 122.195 102.080 122.365 102.250 ;
        RECT 122.555 102.080 122.725 102.250 ;
        RECT 122.915 102.080 123.085 102.250 ;
        RECT 123.275 102.080 123.445 102.250 ;
        RECT 123.635 102.080 123.805 102.250 ;
        RECT 123.995 102.080 124.165 102.250 ;
        RECT 124.600 102.080 124.770 102.250 ;
        RECT 124.960 102.080 125.130 102.250 ;
        RECT 125.320 102.080 125.490 102.250 ;
        RECT 125.680 102.080 125.850 102.250 ;
        RECT 126.040 102.080 126.210 102.250 ;
        RECT 126.400 102.080 126.570 102.250 ;
        RECT 127.165 102.080 127.335 102.250 ;
        RECT 127.525 102.080 127.695 102.250 ;
        RECT 127.885 102.080 128.055 102.250 ;
        RECT 128.245 102.080 128.415 102.250 ;
        RECT 128.605 102.080 128.775 102.250 ;
        RECT 128.965 102.080 129.135 102.250 ;
        RECT 11.020 101.800 11.190 101.970 ;
        RECT 11.705 101.190 41.395 101.720 ;
        RECT 11.100 100.760 11.270 100.930 ;
        RECT 109.770 100.810 109.940 100.980 ;
        RECT 110.130 100.810 110.300 100.980 ;
        RECT 110.490 100.810 110.660 100.980 ;
        RECT 110.850 100.810 111.020 100.980 ;
        RECT 111.210 100.810 111.380 100.980 ;
        RECT 111.570 100.810 111.740 100.980 ;
        RECT 11.100 100.400 11.270 100.570 ;
        RECT 112.175 100.810 112.345 100.980 ;
        RECT 112.535 100.810 112.705 100.980 ;
        RECT 112.895 100.810 113.065 100.980 ;
        RECT 113.255 100.810 113.425 100.980 ;
        RECT 113.615 100.810 113.785 100.980 ;
        RECT 113.975 100.810 114.145 100.980 ;
        RECT 114.740 100.810 114.910 100.980 ;
        RECT 115.100 100.810 115.270 100.980 ;
        RECT 115.460 100.810 115.630 100.980 ;
        RECT 115.820 100.810 115.990 100.980 ;
        RECT 116.180 100.810 116.350 100.980 ;
        RECT 116.540 100.810 116.710 100.980 ;
        RECT 117.145 100.810 117.315 100.980 ;
        RECT 117.505 100.810 117.675 100.980 ;
        RECT 117.865 100.810 118.035 100.980 ;
        RECT 118.225 100.810 118.395 100.980 ;
        RECT 118.585 100.810 118.755 100.980 ;
        RECT 118.945 100.810 119.115 100.980 ;
        RECT 119.710 100.810 119.880 100.980 ;
        RECT 120.070 100.810 120.240 100.980 ;
        RECT 120.430 100.810 120.600 100.980 ;
        RECT 120.790 100.810 120.960 100.980 ;
        RECT 121.150 100.810 121.320 100.980 ;
        RECT 121.510 100.810 121.680 100.980 ;
        RECT 122.115 100.810 122.285 100.980 ;
        RECT 122.475 100.810 122.645 100.980 ;
        RECT 122.835 100.810 123.005 100.980 ;
        RECT 123.195 100.810 123.365 100.980 ;
        RECT 123.555 100.810 123.725 100.980 ;
        RECT 123.915 100.810 124.085 100.980 ;
        RECT 124.680 100.810 124.850 100.980 ;
        RECT 125.040 100.810 125.210 100.980 ;
        RECT 125.400 100.810 125.570 100.980 ;
        RECT 125.760 100.810 125.930 100.980 ;
        RECT 126.120 100.810 126.290 100.980 ;
        RECT 126.480 100.810 126.650 100.980 ;
        RECT 127.085 100.810 127.255 100.980 ;
        RECT 127.445 100.810 127.615 100.980 ;
        RECT 127.805 100.810 127.975 100.980 ;
        RECT 128.165 100.810 128.335 100.980 ;
        RECT 128.525 100.810 128.695 100.980 ;
        RECT 128.885 100.810 129.055 100.980 ;
        RECT 11.100 100.040 11.270 100.210 ;
        RECT 11.100 99.680 11.270 99.850 ;
        RECT 56.250 99.900 56.420 100.070 ;
        RECT 11.100 99.320 11.270 99.490 ;
        RECT 56.935 99.290 86.625 99.820 ;
        RECT 11.705 98.530 41.395 99.060 ;
        RECT 56.330 98.860 56.500 99.030 ;
        RECT 56.330 98.500 56.500 98.670 ;
        RECT 56.330 98.140 56.500 98.310 ;
        RECT 11.665 97.080 51.435 97.970 ;
        RECT 56.330 97.780 56.500 97.950 ;
        RECT 56.330 97.420 56.500 97.590 ;
        RECT 11.100 96.730 11.270 96.900 ;
        RECT 56.935 96.630 86.625 97.160 ;
        RECT 11.100 96.370 11.270 96.540 ;
        RECT 11.100 96.010 11.270 96.180 ;
        RECT 11.100 95.650 11.270 95.820 ;
        RECT 11.100 95.290 11.270 95.460 ;
        RECT 56.895 95.180 96.665 96.070 ;
        RECT 11.100 94.930 11.270 95.100 ;
        RECT 11.100 94.570 11.270 94.740 ;
        RECT 11.100 94.210 11.270 94.380 ;
        RECT 11.100 93.850 11.270 94.020 ;
        RECT 11.100 93.490 11.270 93.660 ;
        RECT 11.100 93.130 11.270 93.300 ;
        RECT 56.330 94.830 56.500 95.000 ;
        RECT 56.330 94.470 56.500 94.640 ;
        RECT 56.330 94.110 56.500 94.280 ;
        RECT 56.330 93.750 56.500 93.920 ;
        RECT 56.330 93.390 56.500 93.560 ;
        RECT 56.330 93.030 56.500 93.200 ;
        RECT 56.330 92.670 56.500 92.840 ;
        RECT 56.330 92.310 56.500 92.480 ;
        RECT 56.330 91.950 56.500 92.120 ;
        RECT 56.330 91.590 56.500 91.760 ;
        RECT 56.330 91.230 56.500 91.400 ;
        RECT 102.625 89.560 102.795 89.730 ;
        RECT 102.985 89.560 103.155 89.730 ;
        RECT 103.345 89.560 103.515 89.730 ;
        RECT 103.705 89.560 103.875 89.730 ;
        RECT 104.065 89.560 104.235 89.730 ;
        RECT 104.425 89.560 104.595 89.730 ;
        RECT 104.785 89.560 104.955 89.730 ;
        RECT 105.145 89.560 105.315 89.730 ;
        RECT 105.505 89.560 105.675 89.730 ;
        RECT 105.865 89.560 106.035 89.730 ;
        RECT 106.225 89.560 106.395 89.730 ;
        RECT 108.815 89.560 108.985 89.730 ;
        RECT 109.175 89.560 109.345 89.730 ;
        RECT 109.535 89.560 109.705 89.730 ;
        RECT 109.895 89.560 110.065 89.730 ;
        RECT 110.255 89.560 110.425 89.730 ;
        RECT 111.295 89.640 111.465 89.810 ;
        RECT 6.630 48.070 7.160 77.760 ;
        RECT 9.290 48.070 9.820 77.760 ;
        RECT 10.380 48.030 11.270 87.800 ;
        RECT 106.575 49.395 107.465 89.165 ;
        RECT 108.025 59.435 108.555 89.125 ;
        RECT 110.685 59.435 111.215 89.125 ;
        RECT 6.380 47.385 6.550 47.555 ;
        RECT 7.420 47.465 7.590 47.635 ;
        RECT 7.780 47.465 7.950 47.635 ;
        RECT 8.140 47.465 8.310 47.635 ;
        RECT 8.500 47.465 8.670 47.635 ;
        RECT 8.860 47.465 9.030 47.635 ;
        RECT 11.450 47.465 11.620 47.635 ;
        RECT 11.810 47.465 11.980 47.635 ;
        RECT 12.170 47.465 12.340 47.635 ;
        RECT 12.530 47.465 12.700 47.635 ;
        RECT 12.890 47.465 13.060 47.635 ;
        RECT 13.250 47.465 13.420 47.635 ;
        RECT 13.610 47.465 13.780 47.635 ;
        RECT 13.970 47.465 14.140 47.635 ;
        RECT 14.330 47.465 14.500 47.635 ;
        RECT 14.690 47.465 14.860 47.635 ;
        RECT 15.050 47.465 15.220 47.635 ;
        RECT 12.680 5.815 13.210 35.505 ;
        RECT 15.340 5.815 15.870 35.505 ;
        RECT 16.430 5.775 17.320 45.545 ;
        RECT 106.575 25.405 106.745 25.575 ;
        RECT 106.575 25.045 106.745 25.215 ;
        RECT 106.575 24.685 106.745 24.855 ;
        RECT 106.575 24.325 106.745 24.495 ;
        RECT 106.575 23.965 106.745 24.135 ;
        RECT 106.575 23.605 106.745 23.775 ;
        RECT 106.575 23.245 106.745 23.415 ;
        RECT 106.575 22.885 106.745 23.055 ;
        RECT 106.575 22.525 106.745 22.695 ;
        RECT 106.575 22.165 106.745 22.335 ;
        RECT 106.575 21.805 106.745 21.975 ;
        RECT 66.410 20.735 106.180 21.625 ;
        RECT 76.450 19.645 106.140 20.175 ;
        RECT 106.575 19.215 106.745 19.385 ;
        RECT 106.575 18.855 106.745 19.025 ;
        RECT 106.575 18.495 106.745 18.665 ;
        RECT 106.575 18.135 106.745 18.305 ;
        RECT 106.575 17.775 106.745 17.945 ;
        RECT 76.450 16.985 106.140 17.515 ;
        RECT 106.655 16.735 106.825 16.905 ;
        RECT 66.360 15.810 66.530 15.980 ;
        RECT 66.360 15.450 66.530 15.620 ;
        RECT 66.360 15.090 66.530 15.260 ;
        RECT 66.360 14.730 66.530 14.900 ;
        RECT 66.360 14.370 66.530 14.540 ;
        RECT 66.360 14.010 66.530 14.180 ;
        RECT 66.360 13.650 66.530 13.820 ;
        RECT 66.360 13.290 66.530 13.460 ;
        RECT 66.360 12.930 66.530 13.100 ;
        RECT 66.360 12.570 66.530 12.740 ;
        RECT 66.360 12.210 66.530 12.380 ;
        RECT 26.195 11.140 65.965 12.030 ;
        RECT 36.235 10.050 65.925 10.580 ;
        RECT 66.360 9.620 66.530 9.790 ;
        RECT 66.360 9.260 66.530 9.430 ;
        RECT 66.360 8.900 66.530 9.070 ;
        RECT 66.360 8.540 66.530 8.710 ;
        RECT 66.360 8.180 66.530 8.350 ;
        RECT 36.235 7.390 65.925 7.920 ;
        RECT 66.440 7.140 66.610 7.310 ;
        RECT 12.430 5.130 12.600 5.300 ;
        RECT 13.470 5.210 13.640 5.380 ;
        RECT 13.830 5.210 14.000 5.380 ;
        RECT 14.190 5.210 14.360 5.380 ;
        RECT 14.550 5.210 14.720 5.380 ;
        RECT 14.910 5.210 15.080 5.380 ;
        RECT 17.500 5.210 17.670 5.380 ;
        RECT 17.860 5.210 18.030 5.380 ;
        RECT 18.220 5.210 18.390 5.380 ;
        RECT 18.580 5.210 18.750 5.380 ;
        RECT 18.940 5.210 19.110 5.380 ;
        RECT 19.300 5.210 19.470 5.380 ;
        RECT 19.660 5.210 19.830 5.380 ;
        RECT 20.020 5.210 20.190 5.380 ;
        RECT 20.380 5.210 20.550 5.380 ;
        RECT 20.740 5.210 20.910 5.380 ;
        RECT 21.100 5.210 21.270 5.380 ;
      LAYER met1 ;
        RECT 9.035 103.885 56.450 106.070 ;
        RECT 102.630 105.455 103.965 105.460 ;
        RECT 102.030 105.090 103.965 105.455 ;
        RECT 102.030 105.085 102.690 105.090 ;
        RECT 2.285 101.700 11.220 103.885 ;
        RECT 2.285 47.585 4.465 101.700 ;
        RECT 11.625 101.160 41.475 101.750 ;
        RECT 6.600 47.990 7.190 77.840 ;
        RECT 9.260 47.950 11.300 100.990 ;
        RECT 54.265 99.800 56.450 103.885 ;
        RECT 56.855 99.260 86.705 99.850 ;
        RECT 11.585 97.050 56.530 99.090 ;
        RECT 103.595 97.190 103.965 105.090 ;
        RECT 55.955 91.170 56.530 97.050 ;
        RECT 56.815 95.150 103.965 97.190 ;
        RECT 109.625 98.770 111.810 103.560 ;
        RECT 112.110 100.770 114.295 104.830 ;
        RECT 114.595 100.770 116.780 106.100 ;
        RECT 117.080 100.770 119.265 107.370 ;
        RECT 119.565 100.770 121.750 107.370 ;
        RECT 122.050 100.770 124.235 106.100 ;
        RECT 139.585 105.005 140.475 105.595 ;
        RECT 124.535 100.770 126.720 104.830 ;
        RECT 127.020 100.770 129.205 103.560 ;
        RECT 136.390 102.450 136.560 102.620 ;
        RECT 109.625 96.585 113.380 98.770 ;
        RECT 102.565 90.105 103.965 95.150 ;
        RECT 111.195 91.795 113.380 96.585 ;
        RECT 102.565 89.530 110.485 90.105 ;
        RECT 111.195 89.610 117.135 91.795 ;
        RECT 2.285 45.400 6.650 47.585 ;
        RECT 7.360 45.625 17.350 47.665 ;
        RECT 4.465 5.330 6.650 45.400 ;
        RECT 12.650 5.735 13.240 35.585 ;
        RECT 15.310 5.695 17.350 45.625 ;
        RECT 66.330 19.615 106.260 21.655 ;
        RECT 26.115 10.020 66.045 12.060 ;
        RECT 26.115 5.410 28.155 10.020 ;
        RECT 66.330 8.120 68.370 19.615 ;
        RECT 106.545 17.715 108.585 89.245 ;
        RECT 110.655 59.355 111.245 89.205 ;
        RECT 76.370 16.955 106.220 17.545 ;
        RECT 114.955 17.005 117.135 89.610 ;
        RECT 106.625 14.820 117.135 17.005 ;
        RECT 36.155 7.360 66.005 7.950 ;
        RECT 106.625 7.410 108.810 14.820 ;
        RECT 4.465 3.145 12.700 5.330 ;
        RECT 13.410 3.910 28.155 5.410 ;
        RECT 66.410 5.225 108.810 7.410 ;
        RECT 66.410 3.145 68.595 5.225 ;
        RECT 10.515 0.965 68.595 3.145 ;
      LAYER met2 ;
        RECT 129.915 100.655 130.115 100.855 ;
        RECT 130.315 100.655 130.515 100.855 ;
        RECT 130.715 100.655 130.915 100.855 ;
        RECT 131.115 100.655 131.315 100.855 ;
        RECT 131.515 100.655 131.715 100.855 ;
        RECT 131.915 100.655 132.115 100.855 ;
        RECT 132.315 100.655 132.515 100.855 ;
        RECT 132.715 100.655 132.915 100.855 ;
        RECT 133.115 100.655 133.315 100.855 ;
        RECT 133.515 100.655 133.715 100.855 ;
        RECT 133.915 100.655 134.115 100.855 ;
        RECT 134.315 100.655 134.515 100.855 ;
        RECT 129.915 100.255 130.115 100.455 ;
        RECT 130.315 100.255 130.515 100.455 ;
        RECT 130.715 100.255 130.915 100.455 ;
        RECT 131.115 100.255 131.315 100.455 ;
        RECT 131.515 100.255 131.715 100.455 ;
        RECT 131.915 100.255 132.115 100.455 ;
        RECT 132.315 100.255 132.515 100.455 ;
        RECT 132.715 100.255 132.915 100.455 ;
        RECT 133.115 100.255 133.315 100.455 ;
        RECT 133.515 100.255 133.715 100.455 ;
        RECT 133.915 100.255 134.115 100.455 ;
        RECT 134.315 100.255 134.515 100.455 ;
  END
END tt_um_wulf_8bit_vco
END LIBRARY

