VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_wulf_8bit_vco
  CLASS BLOCK ;
  FOREIGN tt_um_wulf_8bit_vco ;
  ORIGIN 0.000 0.000 ;
  SIZE 157.320 BY 111.520 ;
  PIN VGND
    ANTENNADIFFAREA 8.540299 ;
    PORT
      LAYER pwell ;
        RECT 11.360 101.910 12.620 103.320 ;
        RECT 11.360 101.810 41.700 101.910 ;
        RECT 11.440 98.330 41.700 101.810 ;
        RECT 56.570 100.010 57.830 101.420 ;
        RECT 56.570 99.910 86.910 100.010 ;
        RECT 56.650 96.430 86.910 99.910 ;
        RECT 110.200 89.390 111.710 89.470 ;
        RECT 106.720 88.210 111.710 89.390 ;
        RECT 6.455 48.980 10.035 78.060 ;
        RECT 106.720 59.130 110.300 88.210 ;
        RECT 5.045 47.800 10.035 48.980 ;
        RECT 5.045 47.720 6.555 47.800 ;
        RECT 12.505 7.880 16.085 36.960 ;
        RECT 75.055 16.890 105.315 20.370 ;
        RECT 75.055 16.790 105.395 16.890 ;
        RECT 104.135 15.380 105.395 16.790 ;
        RECT 11.095 6.700 16.085 7.880 ;
        RECT 34.860 7.295 65.120 10.775 ;
        RECT 34.860 7.195 65.200 7.295 ;
        RECT 11.095 6.620 12.605 6.700 ;
        RECT 63.940 5.785 65.200 7.195 ;
      LAYER li1 ;
        RECT 85.455 106.355 102.475 106.525 ;
        RECT 85.990 105.875 86.160 106.355 ;
        RECT 86.830 105.875 87.000 106.355 ;
        RECT 87.670 105.875 87.840 106.355 ;
        RECT 88.510 105.875 88.680 106.355 ;
        RECT 89.350 105.875 89.520 106.355 ;
        RECT 90.190 105.875 90.360 106.355 ;
        RECT 91.030 105.875 91.200 106.355 ;
        RECT 91.870 105.875 92.040 106.355 ;
        RECT 92.710 105.875 92.880 106.355 ;
        RECT 93.550 105.875 93.720 106.355 ;
        RECT 94.390 105.875 94.560 106.355 ;
        RECT 95.230 105.535 95.400 106.355 ;
        RECT 96.050 105.555 96.380 106.355 ;
        RECT 96.890 105.875 97.220 106.355 ;
        RECT 97.730 105.875 98.060 106.355 ;
        RECT 98.570 105.875 98.900 106.355 ;
        RECT 99.410 105.875 99.740 106.355 ;
        RECT 100.250 105.875 100.580 106.355 ;
        RECT 101.620 105.975 101.950 106.355 ;
        RECT 11.645 102.880 12.335 103.050 ;
        RECT 11.645 102.505 12.335 102.675 ;
        RECT 129.710 101.990 131.890 102.340 ;
        RECT 56.855 100.980 57.545 101.150 ;
        RECT 56.855 100.605 57.545 100.775 ;
        RECT 110.895 88.495 111.065 89.185 ;
        RECT 111.270 88.495 111.440 89.185 ;
        RECT 5.315 48.005 5.485 48.695 ;
        RECT 5.690 48.005 5.860 48.695 ;
        RECT 104.420 16.025 105.110 16.195 ;
        RECT 104.420 15.650 105.110 15.820 ;
        RECT 11.365 6.905 11.535 7.595 ;
        RECT 11.740 6.905 11.910 7.595 ;
        RECT 64.225 6.430 64.915 6.600 ;
        RECT 64.225 6.055 64.915 6.225 ;
      LAYER mcon ;
        RECT 85.600 106.355 85.770 106.525 ;
        RECT 86.060 106.355 86.230 106.525 ;
        RECT 86.520 106.355 86.690 106.525 ;
        RECT 86.980 106.355 87.150 106.525 ;
        RECT 87.440 106.355 87.610 106.525 ;
        RECT 87.900 106.355 88.070 106.525 ;
        RECT 88.360 106.355 88.530 106.525 ;
        RECT 88.820 106.355 88.990 106.525 ;
        RECT 89.280 106.355 89.450 106.525 ;
        RECT 89.740 106.355 89.910 106.525 ;
        RECT 90.200 106.355 90.370 106.525 ;
        RECT 90.660 106.355 90.830 106.525 ;
        RECT 91.120 106.355 91.290 106.525 ;
        RECT 91.580 106.355 91.750 106.525 ;
        RECT 92.040 106.355 92.210 106.525 ;
        RECT 92.500 106.355 92.670 106.525 ;
        RECT 92.960 106.355 93.130 106.525 ;
        RECT 93.420 106.355 93.590 106.525 ;
        RECT 93.880 106.355 94.050 106.525 ;
        RECT 94.340 106.355 94.510 106.525 ;
        RECT 94.800 106.355 94.970 106.525 ;
        RECT 95.260 106.355 95.430 106.525 ;
        RECT 95.720 106.355 95.890 106.525 ;
        RECT 96.180 106.355 96.350 106.525 ;
        RECT 96.640 106.355 96.810 106.525 ;
        RECT 97.100 106.355 97.270 106.525 ;
        RECT 97.560 106.355 97.730 106.525 ;
        RECT 98.020 106.355 98.190 106.525 ;
        RECT 98.480 106.355 98.650 106.525 ;
        RECT 98.940 106.355 99.110 106.525 ;
        RECT 99.400 106.355 99.570 106.525 ;
        RECT 99.860 106.355 100.030 106.525 ;
        RECT 100.320 106.355 100.490 106.525 ;
        RECT 100.780 106.355 100.950 106.525 ;
        RECT 101.240 106.355 101.410 106.525 ;
        RECT 101.700 106.355 101.870 106.525 ;
        RECT 102.160 106.355 102.330 106.525 ;
        RECT 11.725 102.880 11.895 103.050 ;
        RECT 12.085 102.880 12.255 103.050 ;
        RECT 11.725 102.505 11.895 102.675 ;
        RECT 12.085 102.505 12.255 102.675 ;
        RECT 129.820 102.080 129.990 102.250 ;
        RECT 130.180 102.080 130.350 102.250 ;
        RECT 130.540 102.080 130.710 102.250 ;
        RECT 130.900 102.080 131.070 102.250 ;
        RECT 131.260 102.080 131.430 102.250 ;
        RECT 131.620 102.080 131.790 102.250 ;
        RECT 56.935 100.980 57.105 101.150 ;
        RECT 57.295 100.980 57.465 101.150 ;
        RECT 56.935 100.605 57.105 100.775 ;
        RECT 57.295 100.605 57.465 100.775 ;
        RECT 110.895 88.935 111.065 89.105 ;
        RECT 110.895 88.575 111.065 88.745 ;
        RECT 111.270 88.935 111.440 89.105 ;
        RECT 111.270 88.575 111.440 88.745 ;
        RECT 5.315 48.445 5.485 48.615 ;
        RECT 5.315 48.085 5.485 48.255 ;
        RECT 5.690 48.445 5.860 48.615 ;
        RECT 5.690 48.085 5.860 48.255 ;
        RECT 104.500 16.025 104.670 16.195 ;
        RECT 104.860 16.025 105.030 16.195 ;
        RECT 104.500 15.650 104.670 15.820 ;
        RECT 104.860 15.650 105.030 15.820 ;
        RECT 11.365 7.345 11.535 7.515 ;
        RECT 11.365 6.985 11.535 7.155 ;
        RECT 11.740 7.345 11.910 7.515 ;
        RECT 11.740 6.985 11.910 7.155 ;
        RECT 64.305 6.430 64.475 6.600 ;
        RECT 64.665 6.430 64.835 6.600 ;
        RECT 64.305 6.055 64.475 6.225 ;
        RECT 64.665 6.055 64.835 6.225 ;
      LAYER met1 ;
        RECT 43.515 108.930 43.885 109.650 ;
        RECT 46.275 108.930 46.645 109.650 ;
        RECT 49.035 108.930 49.405 109.650 ;
        RECT 51.795 108.930 52.165 109.650 ;
        RECT 54.555 108.930 54.925 109.650 ;
        RECT 57.315 108.930 57.685 109.650 ;
        RECT 60.075 108.930 60.445 109.650 ;
        RECT 62.835 108.930 63.205 109.650 ;
        RECT 65.595 108.930 65.965 109.650 ;
        RECT 68.355 108.930 68.725 109.650 ;
        RECT 71.115 108.930 71.485 109.650 ;
        RECT 73.875 108.930 74.245 109.650 ;
        RECT 76.635 108.930 77.005 109.650 ;
        RECT 79.395 108.930 79.765 109.650 ;
        RECT 82.155 108.930 82.525 109.650 ;
        RECT 85.455 106.200 102.475 106.680 ;
        RECT 11.645 102.475 12.335 103.165 ;
        RECT 129.745 102.005 131.865 102.325 ;
        RECT 56.855 100.575 57.545 101.265 ;
        RECT 110.865 88.495 111.555 89.185 ;
        RECT 5.200 48.005 5.890 48.695 ;
        RECT 104.420 15.535 105.110 16.225 ;
        RECT 11.250 6.905 11.940 7.595 ;
        RECT 64.225 5.940 64.915 6.630 ;
      LAYER via ;
        RECT 43.570 109.335 43.830 109.595 ;
        RECT 43.570 108.985 43.830 109.245 ;
        RECT 46.330 109.335 46.590 109.595 ;
        RECT 46.330 108.985 46.590 109.245 ;
        RECT 49.090 109.335 49.350 109.595 ;
        RECT 49.090 108.985 49.350 109.245 ;
        RECT 51.850 109.335 52.110 109.595 ;
        RECT 51.850 108.985 52.110 109.245 ;
        RECT 54.610 109.335 54.870 109.595 ;
        RECT 54.610 108.985 54.870 109.245 ;
        RECT 57.370 109.335 57.630 109.595 ;
        RECT 57.370 108.985 57.630 109.245 ;
        RECT 60.130 109.335 60.390 109.595 ;
        RECT 60.130 108.985 60.390 109.245 ;
        RECT 62.890 109.335 63.150 109.595 ;
        RECT 62.890 108.985 63.150 109.245 ;
        RECT 65.650 109.335 65.910 109.595 ;
        RECT 65.650 108.985 65.910 109.245 ;
        RECT 68.410 109.335 68.670 109.595 ;
        RECT 68.410 108.985 68.670 109.245 ;
        RECT 71.170 109.335 71.430 109.595 ;
        RECT 71.170 108.985 71.430 109.245 ;
        RECT 73.930 109.335 74.190 109.595 ;
        RECT 73.930 108.985 74.190 109.245 ;
        RECT 76.690 109.335 76.950 109.595 ;
        RECT 76.690 108.985 76.950 109.245 ;
        RECT 79.450 109.335 79.710 109.595 ;
        RECT 79.450 108.985 79.710 109.245 ;
        RECT 82.210 109.335 82.470 109.595 ;
        RECT 82.210 108.985 82.470 109.245 ;
        RECT 85.555 106.310 85.815 106.570 ;
        RECT 86.015 106.310 86.275 106.570 ;
        RECT 86.475 106.310 86.735 106.570 ;
        RECT 86.935 106.310 87.195 106.570 ;
        RECT 87.395 106.310 87.655 106.570 ;
        RECT 87.855 106.310 88.115 106.570 ;
        RECT 88.315 106.310 88.575 106.570 ;
        RECT 88.775 106.310 89.035 106.570 ;
        RECT 89.235 106.310 89.495 106.570 ;
        RECT 89.695 106.310 89.955 106.570 ;
        RECT 90.155 106.310 90.415 106.570 ;
        RECT 90.615 106.310 90.875 106.570 ;
        RECT 91.075 106.310 91.335 106.570 ;
        RECT 91.535 106.310 91.795 106.570 ;
        RECT 91.995 106.310 92.255 106.570 ;
        RECT 92.455 106.310 92.715 106.570 ;
        RECT 92.915 106.310 93.175 106.570 ;
        RECT 93.375 106.310 93.635 106.570 ;
        RECT 93.835 106.310 94.095 106.570 ;
        RECT 94.295 106.310 94.555 106.570 ;
        RECT 94.755 106.310 95.015 106.570 ;
        RECT 95.215 106.310 95.475 106.570 ;
        RECT 95.675 106.310 95.935 106.570 ;
        RECT 96.135 106.310 96.395 106.570 ;
        RECT 96.595 106.310 96.855 106.570 ;
        RECT 97.055 106.310 97.315 106.570 ;
        RECT 97.515 106.310 97.775 106.570 ;
        RECT 97.975 106.310 98.235 106.570 ;
        RECT 98.435 106.310 98.695 106.570 ;
        RECT 98.895 106.310 99.155 106.570 ;
        RECT 99.355 106.310 99.615 106.570 ;
        RECT 99.815 106.310 100.075 106.570 ;
        RECT 100.275 106.310 100.535 106.570 ;
        RECT 100.735 106.310 100.995 106.570 ;
        RECT 101.195 106.310 101.455 106.570 ;
        RECT 101.655 106.310 101.915 106.570 ;
        RECT 102.115 106.310 102.375 106.570 ;
        RECT 11.675 102.875 11.935 103.135 ;
        RECT 12.045 102.875 12.305 103.135 ;
        RECT 11.675 102.505 11.935 102.765 ;
        RECT 12.045 102.505 12.305 102.765 ;
        RECT 129.775 102.035 130.035 102.295 ;
        RECT 130.135 102.035 130.395 102.295 ;
        RECT 130.495 102.035 130.755 102.295 ;
        RECT 130.855 102.035 131.115 102.295 ;
        RECT 131.215 102.035 131.475 102.295 ;
        RECT 131.575 102.035 131.835 102.295 ;
        RECT 56.885 100.975 57.145 101.235 ;
        RECT 57.255 100.975 57.515 101.235 ;
        RECT 56.885 100.605 57.145 100.865 ;
        RECT 57.255 100.605 57.515 100.865 ;
        RECT 110.895 88.895 111.155 89.155 ;
        RECT 111.265 88.895 111.525 89.155 ;
        RECT 110.895 88.525 111.155 88.785 ;
        RECT 111.265 88.525 111.525 88.785 ;
        RECT 5.230 48.405 5.490 48.665 ;
        RECT 5.600 48.405 5.860 48.665 ;
        RECT 5.230 48.035 5.490 48.295 ;
        RECT 5.600 48.035 5.860 48.295 ;
        RECT 104.450 15.935 104.710 16.195 ;
        RECT 104.820 15.935 105.080 16.195 ;
        RECT 104.450 15.565 104.710 15.825 ;
        RECT 104.820 15.565 105.080 15.825 ;
        RECT 11.280 7.305 11.540 7.565 ;
        RECT 11.650 7.305 11.910 7.565 ;
        RECT 11.280 6.935 11.540 7.195 ;
        RECT 11.650 6.935 11.910 7.195 ;
        RECT 64.255 6.340 64.515 6.600 ;
        RECT 64.625 6.340 64.885 6.600 ;
        RECT 64.255 5.970 64.515 6.230 ;
        RECT 64.625 5.970 64.885 6.230 ;
      LAYER met2 ;
        RECT 0.000 106.850 19.320 111.520 ;
        RECT 43.510 106.850 82.530 110.425 ;
        RECT 139.580 106.850 157.320 111.520 ;
        RECT 0.000 105.580 157.320 106.850 ;
        RECT 0.000 101.450 83.460 105.580 ;
        RECT 104.485 104.140 157.320 105.580 ;
        RECT 104.485 101.450 105.130 104.140 ;
        RECT 0.000 100.025 105.130 101.450 ;
        RECT 111.125 100.025 157.320 104.140 ;
        RECT 0.000 93.770 157.320 100.025 ;
        RECT 0.000 89.270 9.595 93.770 ;
        RECT 53.485 91.965 157.320 93.770 ;
        RECT 0.000 46.260 14.520 89.270 ;
        RECT 53.485 88.775 54.850 91.965 ;
        RECT 19.545 86.835 54.850 88.775 ;
        RECT 19.545 48.850 97.000 86.835 ;
        RECT 19.545 46.260 20.610 48.850 ;
        RECT 0.000 5.395 20.610 46.260 ;
        RECT 25.660 47.305 97.000 48.850 ;
        RECT 102.245 47.305 157.320 91.965 ;
        RECT 25.660 29.940 157.320 47.305 ;
        RECT 25.660 24.775 63.180 29.940 ;
        RECT 107.245 24.775 157.320 29.940 ;
        RECT 25.660 20.430 157.320 24.775 ;
        RECT 67.000 15.280 157.320 20.430 ;
        RECT 25.660 5.395 157.320 15.280 ;
        RECT 0.000 0.000 157.320 5.395 ;
      LAYER via2 ;
        RECT 43.560 110.100 43.840 110.380 ;
        RECT 46.320 110.100 46.600 110.380 ;
        RECT 49.080 110.100 49.360 110.380 ;
        RECT 51.840 110.100 52.120 110.380 ;
        RECT 54.600 110.100 54.880 110.380 ;
        RECT 57.360 110.100 57.640 110.380 ;
        RECT 60.120 110.100 60.400 110.380 ;
        RECT 62.880 110.100 63.160 110.380 ;
        RECT 65.640 110.100 65.920 110.380 ;
        RECT 68.400 110.100 68.680 110.380 ;
        RECT 71.160 110.100 71.440 110.380 ;
        RECT 73.920 110.100 74.200 110.380 ;
        RECT 76.680 110.100 76.960 110.380 ;
        RECT 79.440 110.100 79.720 110.380 ;
        RECT 82.200 110.100 82.480 110.380 ;
        RECT 43.560 109.700 43.840 109.980 ;
        RECT 46.320 109.700 46.600 109.980 ;
        RECT 49.080 109.700 49.360 109.980 ;
        RECT 51.840 109.700 52.120 109.980 ;
        RECT 54.600 109.700 54.880 109.980 ;
        RECT 57.360 109.700 57.640 109.980 ;
        RECT 60.120 109.700 60.400 109.980 ;
        RECT 62.880 109.700 63.160 109.980 ;
        RECT 65.640 109.700 65.920 109.980 ;
        RECT 68.400 109.700 68.680 109.980 ;
        RECT 71.160 109.700 71.440 109.980 ;
        RECT 73.920 109.700 74.200 109.980 ;
        RECT 76.680 109.700 76.960 109.980 ;
        RECT 79.440 109.700 79.720 109.980 ;
        RECT 82.200 109.700 82.480 109.980 ;
        RECT 155.580 0.220 157.060 111.300 ;
      LAYER met3 ;
        RECT 43.510 109.650 43.890 111.230 ;
        RECT 46.270 109.650 46.650 111.230 ;
        RECT 49.030 109.650 49.410 111.230 ;
        RECT 51.790 109.650 52.170 111.230 ;
        RECT 54.550 109.650 54.930 111.230 ;
        RECT 57.310 109.650 57.690 111.230 ;
        RECT 60.070 109.650 60.450 111.230 ;
        RECT 62.830 109.650 63.210 111.230 ;
        RECT 65.590 109.650 65.970 111.230 ;
        RECT 68.350 109.650 68.730 111.230 ;
        RECT 71.110 109.650 71.490 111.230 ;
        RECT 73.870 109.650 74.250 111.230 ;
        RECT 76.630 109.650 77.010 111.230 ;
        RECT 79.390 109.650 79.770 111.230 ;
        RECT 82.150 109.650 82.530 111.230 ;
        RECT 155.320 0.000 157.320 111.520 ;
      LAYER via3 ;
        RECT 43.540 110.880 43.860 111.200 ;
        RECT 43.540 110.480 43.860 110.800 ;
        RECT 46.300 110.880 46.620 111.200 ;
        RECT 46.300 110.480 46.620 110.800 ;
        RECT 49.060 110.880 49.380 111.200 ;
        RECT 49.060 110.480 49.380 110.800 ;
        RECT 51.820 110.880 52.140 111.200 ;
        RECT 51.820 110.480 52.140 110.800 ;
        RECT 54.580 110.880 54.900 111.200 ;
        RECT 54.580 110.480 54.900 110.800 ;
        RECT 57.340 110.880 57.660 111.200 ;
        RECT 57.340 110.480 57.660 110.800 ;
        RECT 60.100 110.880 60.420 111.200 ;
        RECT 60.100 110.480 60.420 110.800 ;
        RECT 62.860 110.880 63.180 111.200 ;
        RECT 62.860 110.480 63.180 110.800 ;
        RECT 65.620 110.880 65.940 111.200 ;
        RECT 65.620 110.480 65.940 110.800 ;
        RECT 68.380 110.880 68.700 111.200 ;
        RECT 68.380 110.480 68.700 110.800 ;
        RECT 71.140 110.880 71.460 111.200 ;
        RECT 71.140 110.480 71.460 110.800 ;
        RECT 73.900 110.880 74.220 111.200 ;
        RECT 73.900 110.480 74.220 110.800 ;
        RECT 76.660 110.880 76.980 111.200 ;
        RECT 76.660 110.480 76.980 110.800 ;
        RECT 79.420 110.880 79.740 111.200 ;
        RECT 79.420 110.480 79.740 110.800 ;
        RECT 82.180 110.880 82.500 111.200 ;
        RECT 82.180 110.480 82.500 110.800 ;
        RECT 155.560 0.200 157.080 111.320 ;
      LAYER met4 ;
        RECT 43.550 111.230 43.850 111.520 ;
        RECT 46.310 111.230 46.610 111.520 ;
        RECT 49.070 111.230 49.370 111.520 ;
        RECT 51.830 111.230 52.130 111.520 ;
        RECT 54.590 111.230 54.890 111.520 ;
        RECT 57.350 111.230 57.650 111.520 ;
        RECT 60.110 111.230 60.410 111.520 ;
        RECT 62.870 111.230 63.170 111.520 ;
        RECT 65.630 111.230 65.930 111.520 ;
        RECT 68.390 111.230 68.690 111.520 ;
        RECT 71.150 111.230 71.450 111.520 ;
        RECT 73.910 111.230 74.210 111.520 ;
        RECT 76.670 111.230 76.970 111.520 ;
        RECT 79.430 111.230 79.730 111.520 ;
        RECT 82.190 111.230 82.490 111.520 ;
        RECT 43.510 110.450 43.890 111.230 ;
        RECT 46.270 110.450 46.650 111.230 ;
        RECT 49.030 110.450 49.410 111.230 ;
        RECT 51.790 110.450 52.170 111.230 ;
        RECT 54.550 110.450 54.930 111.230 ;
        RECT 57.310 110.450 57.690 111.230 ;
        RECT 60.070 110.450 60.450 111.230 ;
        RECT 62.830 110.450 63.210 111.230 ;
        RECT 65.590 110.450 65.970 111.230 ;
        RECT 68.350 110.450 68.730 111.230 ;
        RECT 71.110 110.450 71.490 111.230 ;
        RECT 73.870 110.450 74.250 111.230 ;
        RECT 76.630 110.450 77.010 111.230 ;
        RECT 79.390 110.450 79.770 111.230 ;
        RECT 82.150 110.450 82.530 111.230 ;
        RECT 155.320 0.000 157.320 111.520 ;
    END
  END VGND
  PIN clk
    PORT
      LAYER met1 ;
        RECT 134.595 108.930 134.965 109.650 ;
      LAYER via ;
        RECT 134.650 109.335 134.910 109.595 ;
        RECT 134.650 108.985 134.910 109.245 ;
      LAYER met2 ;
        RECT 134.590 108.930 134.970 110.425 ;
      LAYER via2 ;
        RECT 134.640 110.100 134.920 110.380 ;
        RECT 134.640 109.700 134.920 109.980 ;
      LAYER met3 ;
        RECT 134.590 109.650 134.970 111.230 ;
      LAYER via3 ;
        RECT 134.620 110.880 134.940 111.200 ;
        RECT 134.620 110.480 134.940 110.800 ;
      LAYER met4 ;
        RECT 134.630 111.230 134.930 111.520 ;
        RECT 134.590 110.450 134.970 111.230 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met1 ;
        RECT 137.355 108.930 137.725 109.650 ;
      LAYER via ;
        RECT 137.410 109.335 137.670 109.595 ;
        RECT 137.410 108.985 137.670 109.245 ;
      LAYER met2 ;
        RECT 137.350 108.930 137.730 110.425 ;
      LAYER via2 ;
        RECT 137.400 110.100 137.680 110.380 ;
        RECT 137.400 109.700 137.680 109.980 ;
      LAYER met3 ;
        RECT 137.350 109.650 137.730 111.230 ;
      LAYER via3 ;
        RECT 137.380 110.880 137.700 111.200 ;
        RECT 137.380 110.480 137.700 110.800 ;
      LAYER met4 ;
        RECT 137.390 111.230 137.690 111.520 ;
        RECT 137.350 110.450 137.730 111.230 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met1 ;
        RECT 131.835 108.930 132.205 109.650 ;
      LAYER via ;
        RECT 131.890 109.335 132.150 109.595 ;
        RECT 131.890 108.985 132.150 109.245 ;
      LAYER met2 ;
        RECT 131.830 108.930 132.210 110.425 ;
      LAYER via2 ;
        RECT 131.880 110.100 132.160 110.380 ;
        RECT 131.880 109.700 132.160 109.980 ;
      LAYER met3 ;
        RECT 131.830 109.650 132.210 111.230 ;
      LAYER via3 ;
        RECT 131.860 110.880 132.180 111.200 ;
        RECT 131.860 110.480 132.180 110.800 ;
      LAYER met4 ;
        RECT 131.870 111.230 132.170 111.520 ;
        RECT 131.830 110.450 132.210 111.230 ;
    END
  END rst_n
  PIN ui_in[0]
    PORT
      LAYER li1 ;
        RECT 129.710 103.260 131.890 103.610 ;
      LAYER mcon ;
        RECT 129.820 103.350 129.990 103.520 ;
        RECT 130.180 103.350 130.350 103.520 ;
        RECT 130.540 103.350 130.710 103.520 ;
        RECT 130.900 103.350 131.070 103.520 ;
        RECT 131.260 103.350 131.430 103.520 ;
        RECT 131.620 103.350 131.790 103.520 ;
      LAYER met1 ;
        RECT 129.075 108.930 129.445 109.650 ;
        RECT 129.075 108.630 130.055 108.930 ;
        RECT 129.755 103.860 130.055 108.630 ;
        RECT 129.755 103.310 131.860 103.860 ;
      LAYER via ;
        RECT 129.130 109.335 129.390 109.595 ;
        RECT 129.130 108.985 129.390 109.245 ;
      LAYER met2 ;
        RECT 129.070 108.930 129.450 110.425 ;
      LAYER via2 ;
        RECT 129.120 110.100 129.400 110.380 ;
        RECT 129.120 109.700 129.400 109.980 ;
      LAYER met3 ;
        RECT 129.070 109.650 129.450 111.230 ;
      LAYER via3 ;
        RECT 129.100 110.880 129.420 111.200 ;
        RECT 129.100 110.480 129.420 110.800 ;
      LAYER met4 ;
        RECT 129.110 111.230 129.410 111.520 ;
        RECT 129.070 110.450 129.450 111.230 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER li1 ;
        RECT 127.225 104.530 129.405 104.880 ;
      LAYER mcon ;
        RECT 127.335 104.620 127.505 104.790 ;
        RECT 127.695 104.620 127.865 104.790 ;
        RECT 128.055 104.620 128.225 104.790 ;
        RECT 128.415 104.620 128.585 104.790 ;
        RECT 128.775 104.620 128.945 104.790 ;
        RECT 129.135 104.620 129.305 104.790 ;
      LAYER met1 ;
        RECT 126.315 108.930 126.685 109.650 ;
        RECT 126.315 108.630 127.570 108.930 ;
        RECT 127.270 105.130 127.570 108.630 ;
        RECT 127.270 104.580 129.375 105.130 ;
      LAYER via ;
        RECT 126.370 109.335 126.630 109.595 ;
        RECT 126.370 108.985 126.630 109.245 ;
      LAYER met2 ;
        RECT 126.310 108.930 126.690 110.425 ;
      LAYER via2 ;
        RECT 126.360 110.100 126.640 110.380 ;
        RECT 126.360 109.700 126.640 109.980 ;
      LAYER met3 ;
        RECT 126.310 109.650 126.690 111.230 ;
      LAYER via3 ;
        RECT 126.340 110.880 126.660 111.200 ;
        RECT 126.340 110.480 126.660 110.800 ;
      LAYER met4 ;
        RECT 126.350 111.230 126.650 111.520 ;
        RECT 126.310 110.450 126.690 111.230 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER li1 ;
        RECT 124.740 105.800 126.920 106.150 ;
      LAYER mcon ;
        RECT 124.850 105.890 125.020 106.060 ;
        RECT 125.210 105.890 125.380 106.060 ;
        RECT 125.570 105.890 125.740 106.060 ;
        RECT 125.930 105.890 126.100 106.060 ;
        RECT 126.290 105.890 126.460 106.060 ;
        RECT 126.650 105.890 126.820 106.060 ;
      LAYER met1 ;
        RECT 123.555 108.930 123.925 109.650 ;
        RECT 123.555 108.630 125.085 108.930 ;
        RECT 124.785 106.400 125.085 108.630 ;
        RECT 124.785 105.850 126.890 106.400 ;
      LAYER via ;
        RECT 123.610 109.335 123.870 109.595 ;
        RECT 123.610 108.985 123.870 109.245 ;
      LAYER met2 ;
        RECT 123.550 108.930 123.930 110.425 ;
      LAYER via2 ;
        RECT 123.600 110.100 123.880 110.380 ;
        RECT 123.600 109.700 123.880 109.980 ;
      LAYER met3 ;
        RECT 123.550 109.650 123.930 111.230 ;
      LAYER via3 ;
        RECT 123.580 110.880 123.900 111.200 ;
        RECT 123.580 110.480 123.900 110.800 ;
      LAYER met4 ;
        RECT 123.590 111.230 123.890 111.520 ;
        RECT 123.550 110.450 123.930 111.230 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER li1 ;
        RECT 122.255 107.070 124.435 107.420 ;
      LAYER mcon ;
        RECT 122.365 107.160 122.535 107.330 ;
        RECT 122.725 107.160 122.895 107.330 ;
        RECT 123.085 107.160 123.255 107.330 ;
        RECT 123.445 107.160 123.615 107.330 ;
        RECT 123.805 107.160 123.975 107.330 ;
        RECT 124.165 107.160 124.335 107.330 ;
      LAYER met1 ;
        RECT 120.795 108.930 121.165 109.650 ;
        RECT 120.795 108.630 122.600 108.930 ;
        RECT 122.300 107.670 122.600 108.630 ;
        RECT 122.300 107.120 124.405 107.670 ;
      LAYER via ;
        RECT 120.850 109.335 121.110 109.595 ;
        RECT 120.850 108.985 121.110 109.245 ;
      LAYER met2 ;
        RECT 120.790 108.930 121.170 110.425 ;
      LAYER via2 ;
        RECT 120.840 110.100 121.120 110.380 ;
        RECT 120.840 109.700 121.120 109.980 ;
      LAYER met3 ;
        RECT 120.790 109.650 121.170 111.230 ;
      LAYER via3 ;
        RECT 120.820 110.880 121.140 111.200 ;
        RECT 120.820 110.480 121.140 110.800 ;
      LAYER met4 ;
        RECT 120.830 111.230 121.130 111.520 ;
        RECT 120.790 110.450 121.170 111.230 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER li1 ;
        RECT 114.395 107.070 116.575 107.420 ;
      LAYER mcon ;
        RECT 114.490 107.160 114.660 107.330 ;
        RECT 114.850 107.160 115.020 107.330 ;
        RECT 115.210 107.160 115.380 107.330 ;
        RECT 115.570 107.160 115.740 107.330 ;
        RECT 115.930 107.160 116.100 107.330 ;
        RECT 116.290 107.160 116.460 107.330 ;
      LAYER met1 ;
        RECT 118.035 108.930 118.405 109.650 ;
        RECT 116.230 108.630 118.405 108.930 ;
        RECT 116.230 107.670 116.530 108.630 ;
        RECT 114.425 107.120 116.530 107.670 ;
      LAYER via ;
        RECT 118.090 109.335 118.350 109.595 ;
        RECT 118.090 108.985 118.350 109.245 ;
      LAYER met2 ;
        RECT 118.030 108.930 118.410 110.425 ;
      LAYER via2 ;
        RECT 118.080 110.100 118.360 110.380 ;
        RECT 118.080 109.700 118.360 109.980 ;
      LAYER met3 ;
        RECT 118.030 109.650 118.410 111.230 ;
      LAYER via3 ;
        RECT 118.060 110.880 118.380 111.200 ;
        RECT 118.060 110.480 118.380 110.800 ;
      LAYER met4 ;
        RECT 118.070 111.230 118.370 111.520 ;
        RECT 118.030 110.450 118.410 111.230 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER li1 ;
        RECT 111.910 105.800 114.090 106.150 ;
      LAYER mcon ;
        RECT 112.005 105.890 112.175 106.060 ;
        RECT 112.365 105.890 112.535 106.060 ;
        RECT 112.725 105.890 112.895 106.060 ;
        RECT 113.085 105.890 113.255 106.060 ;
        RECT 113.445 105.890 113.615 106.060 ;
        RECT 113.805 105.890 113.975 106.060 ;
      LAYER met1 ;
        RECT 115.275 108.930 115.645 109.650 ;
        RECT 113.745 108.630 115.645 108.930 ;
        RECT 113.745 106.400 114.045 108.630 ;
        RECT 111.940 105.850 114.045 106.400 ;
      LAYER via ;
        RECT 115.330 109.335 115.590 109.595 ;
        RECT 115.330 108.985 115.590 109.245 ;
      LAYER met2 ;
        RECT 115.270 108.930 115.650 110.425 ;
      LAYER via2 ;
        RECT 115.320 110.100 115.600 110.380 ;
        RECT 115.320 109.700 115.600 109.980 ;
      LAYER met3 ;
        RECT 115.270 109.650 115.650 111.230 ;
      LAYER via3 ;
        RECT 115.300 110.880 115.620 111.200 ;
        RECT 115.300 110.480 115.620 110.800 ;
      LAYER met4 ;
        RECT 115.310 111.230 115.610 111.520 ;
        RECT 115.270 110.450 115.650 111.230 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER li1 ;
        RECT 109.425 104.530 111.605 104.880 ;
      LAYER mcon ;
        RECT 109.520 104.620 109.690 104.790 ;
        RECT 109.880 104.620 110.050 104.790 ;
        RECT 110.240 104.620 110.410 104.790 ;
        RECT 110.600 104.620 110.770 104.790 ;
        RECT 110.960 104.620 111.130 104.790 ;
        RECT 111.320 104.620 111.490 104.790 ;
      LAYER met1 ;
        RECT 112.515 108.930 112.885 109.650 ;
        RECT 111.260 108.630 112.885 108.930 ;
        RECT 111.260 105.130 111.560 108.630 ;
        RECT 109.455 104.580 111.560 105.130 ;
      LAYER via ;
        RECT 112.570 109.335 112.830 109.595 ;
        RECT 112.570 108.985 112.830 109.245 ;
      LAYER met2 ;
        RECT 112.510 108.930 112.890 110.425 ;
      LAYER via2 ;
        RECT 112.560 110.100 112.840 110.380 ;
        RECT 112.560 109.700 112.840 109.980 ;
      LAYER met3 ;
        RECT 112.510 109.650 112.890 111.230 ;
      LAYER via3 ;
        RECT 112.540 110.880 112.860 111.200 ;
        RECT 112.540 110.480 112.860 110.800 ;
      LAYER met4 ;
        RECT 112.550 111.230 112.850 111.520 ;
        RECT 112.510 110.450 112.890 111.230 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER li1 ;
        RECT 106.940 103.260 109.120 103.610 ;
      LAYER mcon ;
        RECT 107.035 103.350 107.205 103.520 ;
        RECT 107.395 103.350 107.565 103.520 ;
        RECT 107.755 103.350 107.925 103.520 ;
        RECT 108.115 103.350 108.285 103.520 ;
        RECT 108.475 103.350 108.645 103.520 ;
        RECT 108.835 103.350 109.005 103.520 ;
      LAYER met1 ;
        RECT 109.755 108.930 110.125 109.650 ;
        RECT 108.775 108.630 110.125 108.930 ;
        RECT 108.775 103.860 109.075 108.630 ;
        RECT 106.970 103.310 109.075 103.860 ;
      LAYER via ;
        RECT 109.810 109.335 110.070 109.595 ;
        RECT 109.810 108.985 110.070 109.245 ;
      LAYER met2 ;
        RECT 109.750 108.930 110.130 110.425 ;
      LAYER via2 ;
        RECT 109.800 110.100 110.080 110.380 ;
        RECT 109.800 109.700 110.080 109.980 ;
      LAYER met3 ;
        RECT 109.750 109.650 110.130 111.230 ;
      LAYER via3 ;
        RECT 109.780 110.880 110.100 111.200 ;
        RECT 109.780 110.480 110.100 110.800 ;
      LAYER met4 ;
        RECT 109.790 111.230 110.090 111.520 ;
        RECT 109.750 110.450 110.130 111.230 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met1 ;
        RECT 106.995 108.930 107.365 109.650 ;
      LAYER via ;
        RECT 107.050 109.335 107.310 109.595 ;
        RECT 107.050 108.985 107.310 109.245 ;
      LAYER met2 ;
        RECT 106.990 108.930 107.370 110.425 ;
      LAYER via2 ;
        RECT 107.040 110.100 107.320 110.380 ;
        RECT 107.040 109.700 107.320 109.980 ;
      LAYER met3 ;
        RECT 106.990 109.650 107.370 111.230 ;
      LAYER via3 ;
        RECT 107.020 110.880 107.340 111.200 ;
        RECT 107.020 110.480 107.340 110.800 ;
      LAYER met4 ;
        RECT 107.030 111.230 107.330 111.520 ;
        RECT 106.990 110.450 107.370 111.230 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met1 ;
        RECT 104.235 108.930 104.605 109.650 ;
      LAYER via ;
        RECT 104.290 109.335 104.550 109.595 ;
        RECT 104.290 108.985 104.550 109.245 ;
      LAYER met2 ;
        RECT 104.230 108.930 104.610 110.425 ;
      LAYER via2 ;
        RECT 104.280 110.100 104.560 110.380 ;
        RECT 104.280 109.700 104.560 109.980 ;
      LAYER met3 ;
        RECT 104.230 109.650 104.610 111.230 ;
      LAYER via3 ;
        RECT 104.260 110.880 104.580 111.200 ;
        RECT 104.260 110.480 104.580 110.800 ;
      LAYER met4 ;
        RECT 104.270 111.230 104.570 111.520 ;
        RECT 104.230 110.450 104.610 111.230 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met1 ;
        RECT 101.475 108.930 101.845 109.650 ;
      LAYER via ;
        RECT 101.530 109.335 101.790 109.595 ;
        RECT 101.530 108.985 101.790 109.245 ;
      LAYER met2 ;
        RECT 101.470 108.930 101.850 110.425 ;
      LAYER via2 ;
        RECT 101.520 110.100 101.800 110.380 ;
        RECT 101.520 109.700 101.800 109.980 ;
      LAYER met3 ;
        RECT 101.470 109.650 101.850 111.230 ;
      LAYER via3 ;
        RECT 101.500 110.880 101.820 111.200 ;
        RECT 101.500 110.480 101.820 110.800 ;
      LAYER met4 ;
        RECT 101.510 111.230 101.810 111.520 ;
        RECT 101.470 110.450 101.850 111.230 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met1 ;
        RECT 98.715 108.930 99.085 109.650 ;
      LAYER via ;
        RECT 98.770 109.335 99.030 109.595 ;
        RECT 98.770 108.985 99.030 109.245 ;
      LAYER met2 ;
        RECT 98.710 108.930 99.090 110.425 ;
      LAYER via2 ;
        RECT 98.760 110.100 99.040 110.380 ;
        RECT 98.760 109.700 99.040 109.980 ;
      LAYER met3 ;
        RECT 98.710 109.650 99.090 111.230 ;
      LAYER via3 ;
        RECT 98.740 110.880 99.060 111.200 ;
        RECT 98.740 110.480 99.060 110.800 ;
      LAYER met4 ;
        RECT 98.750 111.230 99.050 111.520 ;
        RECT 98.710 110.450 99.090 111.230 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met1 ;
        RECT 95.955 108.930 96.325 109.650 ;
      LAYER via ;
        RECT 96.010 109.335 96.270 109.595 ;
        RECT 96.010 108.985 96.270 109.245 ;
      LAYER met2 ;
        RECT 95.950 108.930 96.330 110.425 ;
      LAYER via2 ;
        RECT 96.000 110.100 96.280 110.380 ;
        RECT 96.000 109.700 96.280 109.980 ;
      LAYER met3 ;
        RECT 95.950 109.650 96.330 111.230 ;
      LAYER via3 ;
        RECT 95.980 110.880 96.300 111.200 ;
        RECT 95.980 110.480 96.300 110.800 ;
      LAYER met4 ;
        RECT 95.990 111.230 96.290 111.520 ;
        RECT 95.950 110.450 96.330 111.230 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met1 ;
        RECT 93.195 108.930 93.565 109.650 ;
      LAYER via ;
        RECT 93.250 109.335 93.510 109.595 ;
        RECT 93.250 108.985 93.510 109.245 ;
      LAYER met2 ;
        RECT 93.190 108.930 93.570 110.425 ;
      LAYER via2 ;
        RECT 93.240 110.100 93.520 110.380 ;
        RECT 93.240 109.700 93.520 109.980 ;
      LAYER met3 ;
        RECT 93.190 109.650 93.570 111.230 ;
      LAYER via3 ;
        RECT 93.220 110.880 93.540 111.200 ;
        RECT 93.220 110.480 93.540 110.800 ;
      LAYER met4 ;
        RECT 93.230 111.230 93.530 111.520 ;
        RECT 93.190 110.450 93.570 111.230 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met1 ;
        RECT 90.435 108.930 90.805 109.650 ;
      LAYER via ;
        RECT 90.490 109.335 90.750 109.595 ;
        RECT 90.490 108.985 90.750 109.245 ;
      LAYER met2 ;
        RECT 90.430 108.930 90.810 110.425 ;
      LAYER via2 ;
        RECT 90.480 110.100 90.760 110.380 ;
        RECT 90.480 109.700 90.760 109.980 ;
      LAYER met3 ;
        RECT 90.430 109.650 90.810 111.230 ;
      LAYER via3 ;
        RECT 90.460 110.880 90.780 111.200 ;
        RECT 90.460 110.480 90.780 110.800 ;
      LAYER met4 ;
        RECT 90.470 111.230 90.770 111.520 ;
        RECT 90.430 110.450 90.810 111.230 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met1 ;
        RECT 87.675 108.930 88.045 109.650 ;
      LAYER via ;
        RECT 87.730 109.335 87.990 109.595 ;
        RECT 87.730 108.985 87.990 109.245 ;
      LAYER met2 ;
        RECT 87.670 108.930 88.050 110.425 ;
      LAYER via2 ;
        RECT 87.720 110.100 88.000 110.380 ;
        RECT 87.720 109.700 88.000 109.980 ;
      LAYER met3 ;
        RECT 87.670 109.650 88.050 111.230 ;
      LAYER via3 ;
        RECT 87.700 110.880 88.020 111.200 ;
        RECT 87.700 110.480 88.020 110.800 ;
      LAYER met4 ;
        RECT 87.710 111.230 88.010 111.520 ;
        RECT 87.670 110.450 88.050 111.230 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 661.659058 ;
    PORT
      LAYER nwell ;
        RECT 10.850 98.330 11.440 98.335 ;
        RECT 41.700 98.330 51.950 98.335 ;
        RECT 10.850 90.360 51.950 98.330 ;
        RECT 56.060 96.430 56.650 96.435 ;
        RECT 86.910 96.430 97.160 96.435 ;
        RECT 56.060 88.460 97.160 96.430 ;
        RECT 98.750 89.390 106.725 89.980 ;
        RECT 10.030 78.060 18.005 88.310 ;
        RECT 10.035 47.800 18.005 78.060 ;
        RECT 98.750 59.130 106.720 89.390 ;
        RECT 98.750 48.880 106.725 59.130 ;
        RECT 10.030 47.210 18.005 47.800 ;
        RECT 16.080 36.960 24.055 47.210 ;
        RECT 16.085 6.700 24.055 36.960 ;
        RECT 64.805 20.370 105.905 28.340 ;
        RECT 64.805 20.365 75.055 20.370 ;
        RECT 105.315 20.365 105.905 20.370 ;
        RECT 24.610 10.775 65.710 18.745 ;
        RECT 24.610 10.770 34.860 10.775 ;
        RECT 65.120 10.770 65.710 10.775 ;
        RECT 16.080 6.110 24.055 6.700 ;
      LAYER li1 ;
        RECT 85.990 103.805 86.160 104.605 ;
        RECT 86.830 103.805 87.000 104.605 ;
        RECT 87.670 103.805 87.840 104.605 ;
        RECT 88.510 103.805 88.680 104.605 ;
        RECT 89.350 103.805 89.520 104.605 ;
        RECT 90.190 103.805 90.360 104.605 ;
        RECT 91.030 103.805 91.200 104.605 ;
        RECT 91.870 103.805 92.040 104.605 ;
        RECT 92.710 103.805 92.880 104.605 ;
        RECT 93.550 103.805 93.720 104.605 ;
        RECT 94.390 103.805 94.560 104.605 ;
        RECT 95.230 103.805 95.400 104.995 ;
        RECT 96.050 103.805 96.380 104.955 ;
        RECT 96.890 103.805 97.220 104.605 ;
        RECT 97.730 103.805 98.060 104.605 ;
        RECT 98.570 103.805 98.900 104.605 ;
        RECT 99.490 103.805 99.660 104.605 ;
        RECT 100.330 103.805 100.500 104.605 ;
        RECT 101.620 103.805 101.950 104.565 ;
        RECT 85.455 103.635 102.475 103.805 ;
        RECT 107.185 101.985 109.375 102.345 ;
        RECT 11.605 92.055 51.535 92.945 ;
        RECT 11.605 90.880 51.535 91.770 ;
        RECT 56.815 90.155 96.745 91.045 ;
        RECT 56.815 88.980 96.745 89.870 ;
        RECT 15.420 47.965 16.310 87.895 ;
        RECT 16.595 47.965 17.485 87.895 ;
        RECT 99.270 49.295 100.160 89.225 ;
        RECT 100.445 49.295 101.335 89.225 ;
        RECT 21.470 6.865 22.360 46.795 ;
        RECT 22.645 6.865 23.535 46.795 ;
        RECT 65.220 26.930 105.150 27.820 ;
        RECT 65.220 25.755 105.150 26.645 ;
        RECT 25.025 17.335 64.955 18.225 ;
        RECT 25.025 16.160 64.955 17.050 ;
      LAYER mcon ;
        RECT 85.600 103.635 85.770 103.805 ;
        RECT 86.060 103.635 86.230 103.805 ;
        RECT 86.520 103.635 86.690 103.805 ;
        RECT 86.980 103.635 87.150 103.805 ;
        RECT 87.440 103.635 87.610 103.805 ;
        RECT 87.900 103.635 88.070 103.805 ;
        RECT 88.360 103.635 88.530 103.805 ;
        RECT 88.820 103.635 88.990 103.805 ;
        RECT 89.280 103.635 89.450 103.805 ;
        RECT 89.740 103.635 89.910 103.805 ;
        RECT 90.200 103.635 90.370 103.805 ;
        RECT 90.660 103.635 90.830 103.805 ;
        RECT 91.120 103.635 91.290 103.805 ;
        RECT 91.580 103.635 91.750 103.805 ;
        RECT 92.040 103.635 92.210 103.805 ;
        RECT 92.500 103.635 92.670 103.805 ;
        RECT 92.960 103.635 93.130 103.805 ;
        RECT 93.420 103.635 93.590 103.805 ;
        RECT 93.880 103.635 94.050 103.805 ;
        RECT 94.340 103.635 94.510 103.805 ;
        RECT 94.800 103.635 94.970 103.805 ;
        RECT 95.260 103.635 95.430 103.805 ;
        RECT 95.720 103.635 95.890 103.805 ;
        RECT 96.180 103.635 96.350 103.805 ;
        RECT 96.640 103.635 96.810 103.805 ;
        RECT 97.100 103.635 97.270 103.805 ;
        RECT 97.560 103.635 97.730 103.805 ;
        RECT 98.020 103.635 98.190 103.805 ;
        RECT 98.480 103.635 98.650 103.805 ;
        RECT 98.940 103.635 99.110 103.805 ;
        RECT 99.400 103.635 99.570 103.805 ;
        RECT 99.860 103.635 100.030 103.805 ;
        RECT 100.320 103.635 100.490 103.805 ;
        RECT 100.780 103.635 100.950 103.805 ;
        RECT 101.240 103.635 101.410 103.805 ;
        RECT 101.700 103.635 101.870 103.805 ;
        RECT 102.160 103.635 102.330 103.805 ;
        RECT 107.285 102.080 107.455 102.250 ;
        RECT 107.645 102.080 107.815 102.250 ;
        RECT 108.005 102.080 108.175 102.250 ;
        RECT 108.365 102.080 108.535 102.250 ;
        RECT 108.725 102.080 108.895 102.250 ;
        RECT 109.085 102.080 109.255 102.250 ;
        RECT 11.685 92.055 51.455 92.945 ;
        RECT 11.685 90.880 51.455 91.770 ;
        RECT 56.895 90.155 96.665 91.045 ;
        RECT 56.895 88.980 96.665 89.870 ;
        RECT 15.420 48.045 16.310 87.815 ;
        RECT 16.595 48.045 17.485 87.815 ;
        RECT 99.270 49.375 100.160 89.145 ;
        RECT 100.445 49.375 101.335 89.145 ;
        RECT 21.470 6.945 22.360 46.715 ;
        RECT 22.645 6.945 23.535 46.715 ;
        RECT 65.300 26.930 105.070 27.820 ;
        RECT 65.300 25.755 105.070 26.645 ;
        RECT 25.105 17.335 64.875 18.225 ;
        RECT 25.105 16.160 64.875 17.050 ;
      LAYER met1 ;
        RECT 21.435 108.930 21.805 109.650 ;
        RECT 24.195 108.930 24.565 109.650 ;
        RECT 26.955 108.930 27.325 109.650 ;
        RECT 29.715 108.930 30.085 109.650 ;
        RECT 32.475 108.930 32.845 109.650 ;
        RECT 35.235 108.930 35.605 109.650 ;
        RECT 37.995 108.930 38.365 109.650 ;
        RECT 40.755 108.930 41.125 109.650 ;
        RECT 85.455 103.480 102.475 103.960 ;
        RECT 107.210 102.005 109.330 102.325 ;
        RECT 11.625 91.770 51.515 92.975 ;
        RECT 11.605 90.835 51.535 91.770 ;
        RECT 56.835 89.870 96.725 91.075 ;
        RECT 56.815 88.935 96.745 89.870 ;
        RECT 99.225 89.205 100.160 89.225 ;
        RECT 16.595 87.875 17.530 87.895 ;
        RECT 15.390 47.985 17.530 87.875 ;
        RECT 99.225 49.315 101.365 89.205 ;
        RECT 99.225 49.295 100.160 49.315 ;
        RECT 16.595 47.965 17.530 47.985 ;
        RECT 22.645 46.775 23.580 46.795 ;
        RECT 21.440 6.885 23.580 46.775 ;
        RECT 65.220 26.930 105.150 27.865 ;
        RECT 65.240 25.725 105.130 26.930 ;
        RECT 25.025 17.335 64.955 18.270 ;
        RECT 25.045 16.130 64.935 17.335 ;
        RECT 22.645 6.865 23.580 6.885 ;
      LAYER via ;
        RECT 21.490 109.335 21.750 109.595 ;
        RECT 21.490 108.985 21.750 109.245 ;
        RECT 24.250 109.335 24.510 109.595 ;
        RECT 24.250 108.985 24.510 109.245 ;
        RECT 27.010 109.335 27.270 109.595 ;
        RECT 27.010 108.985 27.270 109.245 ;
        RECT 29.770 109.335 30.030 109.595 ;
        RECT 29.770 108.985 30.030 109.245 ;
        RECT 32.530 109.335 32.790 109.595 ;
        RECT 32.530 108.985 32.790 109.245 ;
        RECT 35.290 109.335 35.550 109.595 ;
        RECT 35.290 108.985 35.550 109.245 ;
        RECT 38.050 109.335 38.310 109.595 ;
        RECT 38.050 108.985 38.310 109.245 ;
        RECT 40.810 109.335 41.070 109.595 ;
        RECT 40.810 108.985 41.070 109.245 ;
        RECT 85.555 103.590 85.815 103.850 ;
        RECT 86.015 103.590 86.275 103.850 ;
        RECT 86.475 103.590 86.735 103.850 ;
        RECT 86.935 103.590 87.195 103.850 ;
        RECT 87.395 103.590 87.655 103.850 ;
        RECT 87.855 103.590 88.115 103.850 ;
        RECT 88.315 103.590 88.575 103.850 ;
        RECT 88.775 103.590 89.035 103.850 ;
        RECT 89.235 103.590 89.495 103.850 ;
        RECT 89.695 103.590 89.955 103.850 ;
        RECT 90.155 103.590 90.415 103.850 ;
        RECT 90.615 103.590 90.875 103.850 ;
        RECT 91.075 103.590 91.335 103.850 ;
        RECT 91.535 103.590 91.795 103.850 ;
        RECT 91.995 103.590 92.255 103.850 ;
        RECT 92.455 103.590 92.715 103.850 ;
        RECT 92.915 103.590 93.175 103.850 ;
        RECT 93.375 103.590 93.635 103.850 ;
        RECT 93.835 103.590 94.095 103.850 ;
        RECT 94.295 103.590 94.555 103.850 ;
        RECT 94.755 103.590 95.015 103.850 ;
        RECT 95.215 103.590 95.475 103.850 ;
        RECT 95.675 103.590 95.935 103.850 ;
        RECT 96.135 103.590 96.395 103.850 ;
        RECT 96.595 103.590 96.855 103.850 ;
        RECT 97.055 103.590 97.315 103.850 ;
        RECT 97.515 103.590 97.775 103.850 ;
        RECT 97.975 103.590 98.235 103.850 ;
        RECT 98.435 103.590 98.695 103.850 ;
        RECT 98.895 103.590 99.155 103.850 ;
        RECT 99.355 103.590 99.615 103.850 ;
        RECT 99.815 103.590 100.075 103.850 ;
        RECT 100.275 103.590 100.535 103.850 ;
        RECT 100.735 103.590 100.995 103.850 ;
        RECT 101.195 103.590 101.455 103.850 ;
        RECT 101.655 103.590 101.915 103.850 ;
        RECT 102.115 103.590 102.375 103.850 ;
        RECT 107.240 102.035 107.500 102.295 ;
        RECT 107.600 102.035 107.860 102.295 ;
        RECT 107.960 102.035 108.220 102.295 ;
        RECT 108.320 102.035 108.580 102.295 ;
        RECT 108.680 102.035 108.940 102.295 ;
        RECT 109.040 102.035 109.300 102.295 ;
        RECT 11.640 91.555 11.900 91.815 ;
        RECT 12.000 91.555 12.260 91.815 ;
        RECT 12.360 91.555 12.620 91.815 ;
        RECT 12.720 91.555 12.980 91.815 ;
        RECT 13.080 91.555 13.340 91.815 ;
        RECT 13.440 91.555 13.700 91.815 ;
        RECT 13.800 91.555 14.060 91.815 ;
        RECT 14.160 91.555 14.420 91.815 ;
        RECT 14.520 91.555 14.780 91.815 ;
        RECT 14.880 91.555 15.140 91.815 ;
        RECT 15.240 91.555 15.500 91.815 ;
        RECT 15.600 91.555 15.860 91.815 ;
        RECT 15.960 91.555 16.220 91.815 ;
        RECT 16.320 91.555 16.580 91.815 ;
        RECT 16.680 91.555 16.940 91.815 ;
        RECT 17.040 91.555 17.300 91.815 ;
        RECT 17.400 91.555 17.660 91.815 ;
        RECT 17.760 91.555 18.020 91.815 ;
        RECT 18.120 91.555 18.380 91.815 ;
        RECT 18.480 91.555 18.740 91.815 ;
        RECT 18.840 91.555 19.100 91.815 ;
        RECT 19.200 91.555 19.460 91.815 ;
        RECT 19.560 91.555 19.820 91.815 ;
        RECT 19.920 91.555 20.180 91.815 ;
        RECT 20.280 91.555 20.540 91.815 ;
        RECT 20.640 91.555 20.900 91.815 ;
        RECT 21.000 91.555 21.260 91.815 ;
        RECT 21.360 91.555 21.620 91.815 ;
        RECT 21.720 91.555 21.980 91.815 ;
        RECT 22.080 91.555 22.340 91.815 ;
        RECT 22.440 91.555 22.700 91.815 ;
        RECT 22.800 91.555 23.060 91.815 ;
        RECT 23.160 91.555 23.420 91.815 ;
        RECT 23.520 91.555 23.780 91.815 ;
        RECT 23.880 91.555 24.140 91.815 ;
        RECT 24.240 91.555 24.500 91.815 ;
        RECT 24.600 91.555 24.860 91.815 ;
        RECT 24.960 91.555 25.220 91.815 ;
        RECT 25.320 91.555 25.580 91.815 ;
        RECT 25.680 91.555 25.940 91.815 ;
        RECT 26.040 91.555 26.300 91.815 ;
        RECT 26.400 91.555 26.660 91.815 ;
        RECT 26.760 91.555 27.020 91.815 ;
        RECT 27.120 91.555 27.380 91.815 ;
        RECT 27.480 91.555 27.740 91.815 ;
        RECT 27.840 91.555 28.100 91.815 ;
        RECT 28.200 91.555 28.460 91.815 ;
        RECT 28.560 91.555 28.820 91.815 ;
        RECT 28.920 91.555 29.180 91.815 ;
        RECT 29.280 91.555 29.540 91.815 ;
        RECT 29.640 91.555 29.900 91.815 ;
        RECT 30.000 91.555 30.260 91.815 ;
        RECT 30.360 91.555 30.620 91.815 ;
        RECT 30.720 91.555 30.980 91.815 ;
        RECT 31.080 91.555 31.340 91.815 ;
        RECT 31.440 91.555 31.700 91.815 ;
        RECT 31.800 91.555 32.060 91.815 ;
        RECT 32.160 91.555 32.420 91.815 ;
        RECT 32.520 91.555 32.780 91.815 ;
        RECT 32.880 91.555 33.140 91.815 ;
        RECT 33.240 91.555 33.500 91.815 ;
        RECT 33.600 91.555 33.860 91.815 ;
        RECT 33.960 91.555 34.220 91.815 ;
        RECT 34.320 91.555 34.580 91.815 ;
        RECT 34.680 91.555 34.940 91.815 ;
        RECT 35.040 91.555 35.300 91.815 ;
        RECT 35.400 91.555 35.660 91.815 ;
        RECT 35.760 91.555 36.020 91.815 ;
        RECT 36.120 91.555 36.380 91.815 ;
        RECT 36.480 91.555 36.740 91.815 ;
        RECT 36.840 91.555 37.100 91.815 ;
        RECT 37.200 91.555 37.460 91.815 ;
        RECT 37.560 91.555 37.820 91.815 ;
        RECT 37.920 91.555 38.180 91.815 ;
        RECT 38.280 91.555 38.540 91.815 ;
        RECT 38.640 91.555 38.900 91.815 ;
        RECT 39.000 91.555 39.260 91.815 ;
        RECT 39.360 91.555 39.620 91.815 ;
        RECT 39.720 91.555 39.980 91.815 ;
        RECT 40.080 91.555 40.340 91.815 ;
        RECT 40.440 91.555 40.700 91.815 ;
        RECT 40.800 91.555 41.060 91.815 ;
        RECT 41.160 91.555 41.420 91.815 ;
        RECT 41.520 91.555 41.780 91.815 ;
        RECT 41.880 91.555 42.140 91.815 ;
        RECT 42.240 91.555 42.500 91.815 ;
        RECT 42.600 91.555 42.860 91.815 ;
        RECT 42.960 91.555 43.220 91.815 ;
        RECT 43.320 91.555 43.580 91.815 ;
        RECT 43.680 91.555 43.940 91.815 ;
        RECT 44.040 91.555 44.300 91.815 ;
        RECT 44.400 91.555 44.660 91.815 ;
        RECT 44.760 91.555 45.020 91.815 ;
        RECT 45.120 91.555 45.380 91.815 ;
        RECT 45.480 91.555 45.740 91.815 ;
        RECT 45.840 91.555 46.100 91.815 ;
        RECT 46.200 91.555 46.460 91.815 ;
        RECT 46.560 91.555 46.820 91.815 ;
        RECT 46.920 91.555 47.180 91.815 ;
        RECT 47.280 91.555 47.540 91.815 ;
        RECT 47.640 91.555 47.900 91.815 ;
        RECT 48.000 91.555 48.260 91.815 ;
        RECT 48.360 91.555 48.620 91.815 ;
        RECT 48.720 91.555 48.980 91.815 ;
        RECT 49.080 91.555 49.340 91.815 ;
        RECT 49.440 91.555 49.700 91.815 ;
        RECT 49.800 91.555 50.060 91.815 ;
        RECT 50.160 91.555 50.420 91.815 ;
        RECT 50.520 91.555 50.780 91.815 ;
        RECT 50.880 91.555 51.140 91.815 ;
        RECT 51.240 91.555 51.500 91.815 ;
        RECT 11.640 91.195 11.900 91.455 ;
        RECT 12.000 91.195 12.260 91.455 ;
        RECT 12.360 91.195 12.620 91.455 ;
        RECT 12.720 91.195 12.980 91.455 ;
        RECT 13.080 91.195 13.340 91.455 ;
        RECT 13.440 91.195 13.700 91.455 ;
        RECT 13.800 91.195 14.060 91.455 ;
        RECT 14.160 91.195 14.420 91.455 ;
        RECT 14.520 91.195 14.780 91.455 ;
        RECT 14.880 91.195 15.140 91.455 ;
        RECT 15.240 91.195 15.500 91.455 ;
        RECT 15.600 91.195 15.860 91.455 ;
        RECT 15.960 91.195 16.220 91.455 ;
        RECT 16.320 91.195 16.580 91.455 ;
        RECT 16.680 91.195 16.940 91.455 ;
        RECT 17.040 91.195 17.300 91.455 ;
        RECT 17.400 91.195 17.660 91.455 ;
        RECT 17.760 91.195 18.020 91.455 ;
        RECT 18.120 91.195 18.380 91.455 ;
        RECT 18.480 91.195 18.740 91.455 ;
        RECT 18.840 91.195 19.100 91.455 ;
        RECT 19.200 91.195 19.460 91.455 ;
        RECT 19.560 91.195 19.820 91.455 ;
        RECT 19.920 91.195 20.180 91.455 ;
        RECT 20.280 91.195 20.540 91.455 ;
        RECT 20.640 91.195 20.900 91.455 ;
        RECT 21.000 91.195 21.260 91.455 ;
        RECT 21.360 91.195 21.620 91.455 ;
        RECT 21.720 91.195 21.980 91.455 ;
        RECT 22.080 91.195 22.340 91.455 ;
        RECT 22.440 91.195 22.700 91.455 ;
        RECT 22.800 91.195 23.060 91.455 ;
        RECT 23.160 91.195 23.420 91.455 ;
        RECT 23.520 91.195 23.780 91.455 ;
        RECT 23.880 91.195 24.140 91.455 ;
        RECT 24.240 91.195 24.500 91.455 ;
        RECT 24.600 91.195 24.860 91.455 ;
        RECT 24.960 91.195 25.220 91.455 ;
        RECT 25.320 91.195 25.580 91.455 ;
        RECT 25.680 91.195 25.940 91.455 ;
        RECT 26.040 91.195 26.300 91.455 ;
        RECT 26.400 91.195 26.660 91.455 ;
        RECT 26.760 91.195 27.020 91.455 ;
        RECT 27.120 91.195 27.380 91.455 ;
        RECT 27.480 91.195 27.740 91.455 ;
        RECT 27.840 91.195 28.100 91.455 ;
        RECT 28.200 91.195 28.460 91.455 ;
        RECT 28.560 91.195 28.820 91.455 ;
        RECT 28.920 91.195 29.180 91.455 ;
        RECT 29.280 91.195 29.540 91.455 ;
        RECT 29.640 91.195 29.900 91.455 ;
        RECT 30.000 91.195 30.260 91.455 ;
        RECT 30.360 91.195 30.620 91.455 ;
        RECT 30.720 91.195 30.980 91.455 ;
        RECT 31.080 91.195 31.340 91.455 ;
        RECT 31.440 91.195 31.700 91.455 ;
        RECT 31.800 91.195 32.060 91.455 ;
        RECT 32.160 91.195 32.420 91.455 ;
        RECT 32.520 91.195 32.780 91.455 ;
        RECT 32.880 91.195 33.140 91.455 ;
        RECT 33.240 91.195 33.500 91.455 ;
        RECT 33.600 91.195 33.860 91.455 ;
        RECT 33.960 91.195 34.220 91.455 ;
        RECT 34.320 91.195 34.580 91.455 ;
        RECT 34.680 91.195 34.940 91.455 ;
        RECT 35.040 91.195 35.300 91.455 ;
        RECT 35.400 91.195 35.660 91.455 ;
        RECT 35.760 91.195 36.020 91.455 ;
        RECT 36.120 91.195 36.380 91.455 ;
        RECT 36.480 91.195 36.740 91.455 ;
        RECT 36.840 91.195 37.100 91.455 ;
        RECT 37.200 91.195 37.460 91.455 ;
        RECT 37.560 91.195 37.820 91.455 ;
        RECT 37.920 91.195 38.180 91.455 ;
        RECT 38.280 91.195 38.540 91.455 ;
        RECT 38.640 91.195 38.900 91.455 ;
        RECT 39.000 91.195 39.260 91.455 ;
        RECT 39.360 91.195 39.620 91.455 ;
        RECT 39.720 91.195 39.980 91.455 ;
        RECT 40.080 91.195 40.340 91.455 ;
        RECT 40.440 91.195 40.700 91.455 ;
        RECT 40.800 91.195 41.060 91.455 ;
        RECT 41.160 91.195 41.420 91.455 ;
        RECT 41.520 91.195 41.780 91.455 ;
        RECT 41.880 91.195 42.140 91.455 ;
        RECT 42.240 91.195 42.500 91.455 ;
        RECT 42.600 91.195 42.860 91.455 ;
        RECT 42.960 91.195 43.220 91.455 ;
        RECT 43.320 91.195 43.580 91.455 ;
        RECT 43.680 91.195 43.940 91.455 ;
        RECT 44.040 91.195 44.300 91.455 ;
        RECT 44.400 91.195 44.660 91.455 ;
        RECT 44.760 91.195 45.020 91.455 ;
        RECT 45.120 91.195 45.380 91.455 ;
        RECT 45.480 91.195 45.740 91.455 ;
        RECT 45.840 91.195 46.100 91.455 ;
        RECT 46.200 91.195 46.460 91.455 ;
        RECT 46.560 91.195 46.820 91.455 ;
        RECT 46.920 91.195 47.180 91.455 ;
        RECT 47.280 91.195 47.540 91.455 ;
        RECT 47.640 91.195 47.900 91.455 ;
        RECT 48.000 91.195 48.260 91.455 ;
        RECT 48.360 91.195 48.620 91.455 ;
        RECT 48.720 91.195 48.980 91.455 ;
        RECT 49.080 91.195 49.340 91.455 ;
        RECT 49.440 91.195 49.700 91.455 ;
        RECT 49.800 91.195 50.060 91.455 ;
        RECT 50.160 91.195 50.420 91.455 ;
        RECT 50.520 91.195 50.780 91.455 ;
        RECT 50.880 91.195 51.140 91.455 ;
        RECT 51.240 91.195 51.500 91.455 ;
        RECT 11.640 90.835 11.900 91.095 ;
        RECT 12.000 90.835 12.260 91.095 ;
        RECT 12.360 90.835 12.620 91.095 ;
        RECT 12.720 90.835 12.980 91.095 ;
        RECT 13.080 90.835 13.340 91.095 ;
        RECT 13.440 90.835 13.700 91.095 ;
        RECT 13.800 90.835 14.060 91.095 ;
        RECT 14.160 90.835 14.420 91.095 ;
        RECT 14.520 90.835 14.780 91.095 ;
        RECT 14.880 90.835 15.140 91.095 ;
        RECT 15.240 90.835 15.500 91.095 ;
        RECT 15.600 90.835 15.860 91.095 ;
        RECT 15.960 90.835 16.220 91.095 ;
        RECT 16.320 90.835 16.580 91.095 ;
        RECT 16.680 90.835 16.940 91.095 ;
        RECT 17.040 90.835 17.300 91.095 ;
        RECT 17.400 90.835 17.660 91.095 ;
        RECT 17.760 90.835 18.020 91.095 ;
        RECT 18.120 90.835 18.380 91.095 ;
        RECT 18.480 90.835 18.740 91.095 ;
        RECT 18.840 90.835 19.100 91.095 ;
        RECT 19.200 90.835 19.460 91.095 ;
        RECT 19.560 90.835 19.820 91.095 ;
        RECT 19.920 90.835 20.180 91.095 ;
        RECT 20.280 90.835 20.540 91.095 ;
        RECT 20.640 90.835 20.900 91.095 ;
        RECT 21.000 90.835 21.260 91.095 ;
        RECT 21.360 90.835 21.620 91.095 ;
        RECT 21.720 90.835 21.980 91.095 ;
        RECT 22.080 90.835 22.340 91.095 ;
        RECT 22.440 90.835 22.700 91.095 ;
        RECT 22.800 90.835 23.060 91.095 ;
        RECT 23.160 90.835 23.420 91.095 ;
        RECT 23.520 90.835 23.780 91.095 ;
        RECT 23.880 90.835 24.140 91.095 ;
        RECT 24.240 90.835 24.500 91.095 ;
        RECT 24.600 90.835 24.860 91.095 ;
        RECT 24.960 90.835 25.220 91.095 ;
        RECT 25.320 90.835 25.580 91.095 ;
        RECT 25.680 90.835 25.940 91.095 ;
        RECT 26.040 90.835 26.300 91.095 ;
        RECT 26.400 90.835 26.660 91.095 ;
        RECT 26.760 90.835 27.020 91.095 ;
        RECT 27.120 90.835 27.380 91.095 ;
        RECT 27.480 90.835 27.740 91.095 ;
        RECT 27.840 90.835 28.100 91.095 ;
        RECT 28.200 90.835 28.460 91.095 ;
        RECT 28.560 90.835 28.820 91.095 ;
        RECT 28.920 90.835 29.180 91.095 ;
        RECT 29.280 90.835 29.540 91.095 ;
        RECT 29.640 90.835 29.900 91.095 ;
        RECT 30.000 90.835 30.260 91.095 ;
        RECT 30.360 90.835 30.620 91.095 ;
        RECT 30.720 90.835 30.980 91.095 ;
        RECT 31.080 90.835 31.340 91.095 ;
        RECT 31.440 90.835 31.700 91.095 ;
        RECT 31.800 90.835 32.060 91.095 ;
        RECT 32.160 90.835 32.420 91.095 ;
        RECT 32.520 90.835 32.780 91.095 ;
        RECT 32.880 90.835 33.140 91.095 ;
        RECT 33.240 90.835 33.500 91.095 ;
        RECT 33.600 90.835 33.860 91.095 ;
        RECT 33.960 90.835 34.220 91.095 ;
        RECT 34.320 90.835 34.580 91.095 ;
        RECT 34.680 90.835 34.940 91.095 ;
        RECT 35.040 90.835 35.300 91.095 ;
        RECT 35.400 90.835 35.660 91.095 ;
        RECT 35.760 90.835 36.020 91.095 ;
        RECT 36.120 90.835 36.380 91.095 ;
        RECT 36.480 90.835 36.740 91.095 ;
        RECT 36.840 90.835 37.100 91.095 ;
        RECT 37.200 90.835 37.460 91.095 ;
        RECT 37.560 90.835 37.820 91.095 ;
        RECT 37.920 90.835 38.180 91.095 ;
        RECT 38.280 90.835 38.540 91.095 ;
        RECT 38.640 90.835 38.900 91.095 ;
        RECT 39.000 90.835 39.260 91.095 ;
        RECT 39.360 90.835 39.620 91.095 ;
        RECT 39.720 90.835 39.980 91.095 ;
        RECT 40.080 90.835 40.340 91.095 ;
        RECT 40.440 90.835 40.700 91.095 ;
        RECT 40.800 90.835 41.060 91.095 ;
        RECT 41.160 90.835 41.420 91.095 ;
        RECT 41.520 90.835 41.780 91.095 ;
        RECT 41.880 90.835 42.140 91.095 ;
        RECT 42.240 90.835 42.500 91.095 ;
        RECT 42.600 90.835 42.860 91.095 ;
        RECT 42.960 90.835 43.220 91.095 ;
        RECT 43.320 90.835 43.580 91.095 ;
        RECT 43.680 90.835 43.940 91.095 ;
        RECT 44.040 90.835 44.300 91.095 ;
        RECT 44.400 90.835 44.660 91.095 ;
        RECT 44.760 90.835 45.020 91.095 ;
        RECT 45.120 90.835 45.380 91.095 ;
        RECT 45.480 90.835 45.740 91.095 ;
        RECT 45.840 90.835 46.100 91.095 ;
        RECT 46.200 90.835 46.460 91.095 ;
        RECT 46.560 90.835 46.820 91.095 ;
        RECT 46.920 90.835 47.180 91.095 ;
        RECT 47.280 90.835 47.540 91.095 ;
        RECT 47.640 90.835 47.900 91.095 ;
        RECT 48.000 90.835 48.260 91.095 ;
        RECT 48.360 90.835 48.620 91.095 ;
        RECT 48.720 90.835 48.980 91.095 ;
        RECT 49.080 90.835 49.340 91.095 ;
        RECT 49.440 90.835 49.700 91.095 ;
        RECT 49.800 90.835 50.060 91.095 ;
        RECT 50.160 90.835 50.420 91.095 ;
        RECT 50.520 90.835 50.780 91.095 ;
        RECT 50.880 90.835 51.140 91.095 ;
        RECT 51.240 90.835 51.500 91.095 ;
        RECT 56.850 89.655 57.110 89.915 ;
        RECT 57.210 89.655 57.470 89.915 ;
        RECT 57.570 89.655 57.830 89.915 ;
        RECT 57.930 89.655 58.190 89.915 ;
        RECT 58.290 89.655 58.550 89.915 ;
        RECT 58.650 89.655 58.910 89.915 ;
        RECT 59.010 89.655 59.270 89.915 ;
        RECT 59.370 89.655 59.630 89.915 ;
        RECT 59.730 89.655 59.990 89.915 ;
        RECT 60.090 89.655 60.350 89.915 ;
        RECT 60.450 89.655 60.710 89.915 ;
        RECT 60.810 89.655 61.070 89.915 ;
        RECT 61.170 89.655 61.430 89.915 ;
        RECT 61.530 89.655 61.790 89.915 ;
        RECT 61.890 89.655 62.150 89.915 ;
        RECT 62.250 89.655 62.510 89.915 ;
        RECT 62.610 89.655 62.870 89.915 ;
        RECT 62.970 89.655 63.230 89.915 ;
        RECT 63.330 89.655 63.590 89.915 ;
        RECT 63.690 89.655 63.950 89.915 ;
        RECT 64.050 89.655 64.310 89.915 ;
        RECT 64.410 89.655 64.670 89.915 ;
        RECT 64.770 89.655 65.030 89.915 ;
        RECT 65.130 89.655 65.390 89.915 ;
        RECT 65.490 89.655 65.750 89.915 ;
        RECT 65.850 89.655 66.110 89.915 ;
        RECT 66.210 89.655 66.470 89.915 ;
        RECT 66.570 89.655 66.830 89.915 ;
        RECT 66.930 89.655 67.190 89.915 ;
        RECT 67.290 89.655 67.550 89.915 ;
        RECT 67.650 89.655 67.910 89.915 ;
        RECT 68.010 89.655 68.270 89.915 ;
        RECT 68.370 89.655 68.630 89.915 ;
        RECT 68.730 89.655 68.990 89.915 ;
        RECT 69.090 89.655 69.350 89.915 ;
        RECT 69.450 89.655 69.710 89.915 ;
        RECT 69.810 89.655 70.070 89.915 ;
        RECT 70.170 89.655 70.430 89.915 ;
        RECT 70.530 89.655 70.790 89.915 ;
        RECT 70.890 89.655 71.150 89.915 ;
        RECT 71.250 89.655 71.510 89.915 ;
        RECT 71.610 89.655 71.870 89.915 ;
        RECT 71.970 89.655 72.230 89.915 ;
        RECT 72.330 89.655 72.590 89.915 ;
        RECT 72.690 89.655 72.950 89.915 ;
        RECT 73.050 89.655 73.310 89.915 ;
        RECT 73.410 89.655 73.670 89.915 ;
        RECT 73.770 89.655 74.030 89.915 ;
        RECT 74.130 89.655 74.390 89.915 ;
        RECT 74.490 89.655 74.750 89.915 ;
        RECT 74.850 89.655 75.110 89.915 ;
        RECT 75.210 89.655 75.470 89.915 ;
        RECT 75.570 89.655 75.830 89.915 ;
        RECT 75.930 89.655 76.190 89.915 ;
        RECT 76.290 89.655 76.550 89.915 ;
        RECT 76.650 89.655 76.910 89.915 ;
        RECT 77.010 89.655 77.270 89.915 ;
        RECT 77.370 89.655 77.630 89.915 ;
        RECT 77.730 89.655 77.990 89.915 ;
        RECT 78.090 89.655 78.350 89.915 ;
        RECT 78.450 89.655 78.710 89.915 ;
        RECT 78.810 89.655 79.070 89.915 ;
        RECT 79.170 89.655 79.430 89.915 ;
        RECT 79.530 89.655 79.790 89.915 ;
        RECT 79.890 89.655 80.150 89.915 ;
        RECT 80.250 89.655 80.510 89.915 ;
        RECT 80.610 89.655 80.870 89.915 ;
        RECT 80.970 89.655 81.230 89.915 ;
        RECT 81.330 89.655 81.590 89.915 ;
        RECT 81.690 89.655 81.950 89.915 ;
        RECT 82.050 89.655 82.310 89.915 ;
        RECT 82.410 89.655 82.670 89.915 ;
        RECT 82.770 89.655 83.030 89.915 ;
        RECT 83.130 89.655 83.390 89.915 ;
        RECT 83.490 89.655 83.750 89.915 ;
        RECT 83.850 89.655 84.110 89.915 ;
        RECT 84.210 89.655 84.470 89.915 ;
        RECT 84.570 89.655 84.830 89.915 ;
        RECT 84.930 89.655 85.190 89.915 ;
        RECT 85.290 89.655 85.550 89.915 ;
        RECT 85.650 89.655 85.910 89.915 ;
        RECT 86.010 89.655 86.270 89.915 ;
        RECT 86.370 89.655 86.630 89.915 ;
        RECT 86.730 89.655 86.990 89.915 ;
        RECT 87.090 89.655 87.350 89.915 ;
        RECT 87.450 89.655 87.710 89.915 ;
        RECT 87.810 89.655 88.070 89.915 ;
        RECT 88.170 89.655 88.430 89.915 ;
        RECT 88.530 89.655 88.790 89.915 ;
        RECT 88.890 89.655 89.150 89.915 ;
        RECT 89.250 89.655 89.510 89.915 ;
        RECT 89.610 89.655 89.870 89.915 ;
        RECT 89.970 89.655 90.230 89.915 ;
        RECT 90.330 89.655 90.590 89.915 ;
        RECT 90.690 89.655 90.950 89.915 ;
        RECT 91.050 89.655 91.310 89.915 ;
        RECT 91.410 89.655 91.670 89.915 ;
        RECT 91.770 89.655 92.030 89.915 ;
        RECT 92.130 89.655 92.390 89.915 ;
        RECT 92.490 89.655 92.750 89.915 ;
        RECT 92.850 89.655 93.110 89.915 ;
        RECT 93.210 89.655 93.470 89.915 ;
        RECT 93.570 89.655 93.830 89.915 ;
        RECT 93.930 89.655 94.190 89.915 ;
        RECT 94.290 89.655 94.550 89.915 ;
        RECT 94.650 89.655 94.910 89.915 ;
        RECT 95.010 89.655 95.270 89.915 ;
        RECT 95.370 89.655 95.630 89.915 ;
        RECT 95.730 89.655 95.990 89.915 ;
        RECT 96.090 89.655 96.350 89.915 ;
        RECT 96.450 89.655 96.710 89.915 ;
        RECT 56.850 89.295 57.110 89.555 ;
        RECT 57.210 89.295 57.470 89.555 ;
        RECT 57.570 89.295 57.830 89.555 ;
        RECT 57.930 89.295 58.190 89.555 ;
        RECT 58.290 89.295 58.550 89.555 ;
        RECT 58.650 89.295 58.910 89.555 ;
        RECT 59.010 89.295 59.270 89.555 ;
        RECT 59.370 89.295 59.630 89.555 ;
        RECT 59.730 89.295 59.990 89.555 ;
        RECT 60.090 89.295 60.350 89.555 ;
        RECT 60.450 89.295 60.710 89.555 ;
        RECT 60.810 89.295 61.070 89.555 ;
        RECT 61.170 89.295 61.430 89.555 ;
        RECT 61.530 89.295 61.790 89.555 ;
        RECT 61.890 89.295 62.150 89.555 ;
        RECT 62.250 89.295 62.510 89.555 ;
        RECT 62.610 89.295 62.870 89.555 ;
        RECT 62.970 89.295 63.230 89.555 ;
        RECT 63.330 89.295 63.590 89.555 ;
        RECT 63.690 89.295 63.950 89.555 ;
        RECT 64.050 89.295 64.310 89.555 ;
        RECT 64.410 89.295 64.670 89.555 ;
        RECT 64.770 89.295 65.030 89.555 ;
        RECT 65.130 89.295 65.390 89.555 ;
        RECT 65.490 89.295 65.750 89.555 ;
        RECT 65.850 89.295 66.110 89.555 ;
        RECT 66.210 89.295 66.470 89.555 ;
        RECT 66.570 89.295 66.830 89.555 ;
        RECT 66.930 89.295 67.190 89.555 ;
        RECT 67.290 89.295 67.550 89.555 ;
        RECT 67.650 89.295 67.910 89.555 ;
        RECT 68.010 89.295 68.270 89.555 ;
        RECT 68.370 89.295 68.630 89.555 ;
        RECT 68.730 89.295 68.990 89.555 ;
        RECT 69.090 89.295 69.350 89.555 ;
        RECT 69.450 89.295 69.710 89.555 ;
        RECT 69.810 89.295 70.070 89.555 ;
        RECT 70.170 89.295 70.430 89.555 ;
        RECT 70.530 89.295 70.790 89.555 ;
        RECT 70.890 89.295 71.150 89.555 ;
        RECT 71.250 89.295 71.510 89.555 ;
        RECT 71.610 89.295 71.870 89.555 ;
        RECT 71.970 89.295 72.230 89.555 ;
        RECT 72.330 89.295 72.590 89.555 ;
        RECT 72.690 89.295 72.950 89.555 ;
        RECT 73.050 89.295 73.310 89.555 ;
        RECT 73.410 89.295 73.670 89.555 ;
        RECT 73.770 89.295 74.030 89.555 ;
        RECT 74.130 89.295 74.390 89.555 ;
        RECT 74.490 89.295 74.750 89.555 ;
        RECT 74.850 89.295 75.110 89.555 ;
        RECT 75.210 89.295 75.470 89.555 ;
        RECT 75.570 89.295 75.830 89.555 ;
        RECT 75.930 89.295 76.190 89.555 ;
        RECT 76.290 89.295 76.550 89.555 ;
        RECT 76.650 89.295 76.910 89.555 ;
        RECT 77.010 89.295 77.270 89.555 ;
        RECT 77.370 89.295 77.630 89.555 ;
        RECT 77.730 89.295 77.990 89.555 ;
        RECT 78.090 89.295 78.350 89.555 ;
        RECT 78.450 89.295 78.710 89.555 ;
        RECT 78.810 89.295 79.070 89.555 ;
        RECT 79.170 89.295 79.430 89.555 ;
        RECT 79.530 89.295 79.790 89.555 ;
        RECT 79.890 89.295 80.150 89.555 ;
        RECT 80.250 89.295 80.510 89.555 ;
        RECT 80.610 89.295 80.870 89.555 ;
        RECT 80.970 89.295 81.230 89.555 ;
        RECT 81.330 89.295 81.590 89.555 ;
        RECT 81.690 89.295 81.950 89.555 ;
        RECT 82.050 89.295 82.310 89.555 ;
        RECT 82.410 89.295 82.670 89.555 ;
        RECT 82.770 89.295 83.030 89.555 ;
        RECT 83.130 89.295 83.390 89.555 ;
        RECT 83.490 89.295 83.750 89.555 ;
        RECT 83.850 89.295 84.110 89.555 ;
        RECT 84.210 89.295 84.470 89.555 ;
        RECT 84.570 89.295 84.830 89.555 ;
        RECT 84.930 89.295 85.190 89.555 ;
        RECT 85.290 89.295 85.550 89.555 ;
        RECT 85.650 89.295 85.910 89.555 ;
        RECT 86.010 89.295 86.270 89.555 ;
        RECT 86.370 89.295 86.630 89.555 ;
        RECT 86.730 89.295 86.990 89.555 ;
        RECT 87.090 89.295 87.350 89.555 ;
        RECT 87.450 89.295 87.710 89.555 ;
        RECT 87.810 89.295 88.070 89.555 ;
        RECT 88.170 89.295 88.430 89.555 ;
        RECT 88.530 89.295 88.790 89.555 ;
        RECT 88.890 89.295 89.150 89.555 ;
        RECT 89.250 89.295 89.510 89.555 ;
        RECT 89.610 89.295 89.870 89.555 ;
        RECT 89.970 89.295 90.230 89.555 ;
        RECT 90.330 89.295 90.590 89.555 ;
        RECT 90.690 89.295 90.950 89.555 ;
        RECT 91.050 89.295 91.310 89.555 ;
        RECT 91.410 89.295 91.670 89.555 ;
        RECT 91.770 89.295 92.030 89.555 ;
        RECT 92.130 89.295 92.390 89.555 ;
        RECT 92.490 89.295 92.750 89.555 ;
        RECT 92.850 89.295 93.110 89.555 ;
        RECT 93.210 89.295 93.470 89.555 ;
        RECT 93.570 89.295 93.830 89.555 ;
        RECT 93.930 89.295 94.190 89.555 ;
        RECT 94.290 89.295 94.550 89.555 ;
        RECT 94.650 89.295 94.910 89.555 ;
        RECT 95.010 89.295 95.270 89.555 ;
        RECT 95.370 89.295 95.630 89.555 ;
        RECT 95.730 89.295 95.990 89.555 ;
        RECT 96.090 89.295 96.350 89.555 ;
        RECT 96.450 89.295 96.710 89.555 ;
        RECT 56.850 88.935 57.110 89.195 ;
        RECT 57.210 88.935 57.470 89.195 ;
        RECT 57.570 88.935 57.830 89.195 ;
        RECT 57.930 88.935 58.190 89.195 ;
        RECT 58.290 88.935 58.550 89.195 ;
        RECT 58.650 88.935 58.910 89.195 ;
        RECT 59.010 88.935 59.270 89.195 ;
        RECT 59.370 88.935 59.630 89.195 ;
        RECT 59.730 88.935 59.990 89.195 ;
        RECT 60.090 88.935 60.350 89.195 ;
        RECT 60.450 88.935 60.710 89.195 ;
        RECT 60.810 88.935 61.070 89.195 ;
        RECT 61.170 88.935 61.430 89.195 ;
        RECT 61.530 88.935 61.790 89.195 ;
        RECT 61.890 88.935 62.150 89.195 ;
        RECT 62.250 88.935 62.510 89.195 ;
        RECT 62.610 88.935 62.870 89.195 ;
        RECT 62.970 88.935 63.230 89.195 ;
        RECT 63.330 88.935 63.590 89.195 ;
        RECT 63.690 88.935 63.950 89.195 ;
        RECT 64.050 88.935 64.310 89.195 ;
        RECT 64.410 88.935 64.670 89.195 ;
        RECT 64.770 88.935 65.030 89.195 ;
        RECT 65.130 88.935 65.390 89.195 ;
        RECT 65.490 88.935 65.750 89.195 ;
        RECT 65.850 88.935 66.110 89.195 ;
        RECT 66.210 88.935 66.470 89.195 ;
        RECT 66.570 88.935 66.830 89.195 ;
        RECT 66.930 88.935 67.190 89.195 ;
        RECT 67.290 88.935 67.550 89.195 ;
        RECT 67.650 88.935 67.910 89.195 ;
        RECT 68.010 88.935 68.270 89.195 ;
        RECT 68.370 88.935 68.630 89.195 ;
        RECT 68.730 88.935 68.990 89.195 ;
        RECT 69.090 88.935 69.350 89.195 ;
        RECT 69.450 88.935 69.710 89.195 ;
        RECT 69.810 88.935 70.070 89.195 ;
        RECT 70.170 88.935 70.430 89.195 ;
        RECT 70.530 88.935 70.790 89.195 ;
        RECT 70.890 88.935 71.150 89.195 ;
        RECT 71.250 88.935 71.510 89.195 ;
        RECT 71.610 88.935 71.870 89.195 ;
        RECT 71.970 88.935 72.230 89.195 ;
        RECT 72.330 88.935 72.590 89.195 ;
        RECT 72.690 88.935 72.950 89.195 ;
        RECT 73.050 88.935 73.310 89.195 ;
        RECT 73.410 88.935 73.670 89.195 ;
        RECT 73.770 88.935 74.030 89.195 ;
        RECT 74.130 88.935 74.390 89.195 ;
        RECT 74.490 88.935 74.750 89.195 ;
        RECT 74.850 88.935 75.110 89.195 ;
        RECT 75.210 88.935 75.470 89.195 ;
        RECT 75.570 88.935 75.830 89.195 ;
        RECT 75.930 88.935 76.190 89.195 ;
        RECT 76.290 88.935 76.550 89.195 ;
        RECT 76.650 88.935 76.910 89.195 ;
        RECT 77.010 88.935 77.270 89.195 ;
        RECT 77.370 88.935 77.630 89.195 ;
        RECT 77.730 88.935 77.990 89.195 ;
        RECT 78.090 88.935 78.350 89.195 ;
        RECT 78.450 88.935 78.710 89.195 ;
        RECT 78.810 88.935 79.070 89.195 ;
        RECT 79.170 88.935 79.430 89.195 ;
        RECT 79.530 88.935 79.790 89.195 ;
        RECT 79.890 88.935 80.150 89.195 ;
        RECT 80.250 88.935 80.510 89.195 ;
        RECT 80.610 88.935 80.870 89.195 ;
        RECT 80.970 88.935 81.230 89.195 ;
        RECT 81.330 88.935 81.590 89.195 ;
        RECT 81.690 88.935 81.950 89.195 ;
        RECT 82.050 88.935 82.310 89.195 ;
        RECT 82.410 88.935 82.670 89.195 ;
        RECT 82.770 88.935 83.030 89.195 ;
        RECT 83.130 88.935 83.390 89.195 ;
        RECT 83.490 88.935 83.750 89.195 ;
        RECT 83.850 88.935 84.110 89.195 ;
        RECT 84.210 88.935 84.470 89.195 ;
        RECT 84.570 88.935 84.830 89.195 ;
        RECT 84.930 88.935 85.190 89.195 ;
        RECT 85.290 88.935 85.550 89.195 ;
        RECT 85.650 88.935 85.910 89.195 ;
        RECT 86.010 88.935 86.270 89.195 ;
        RECT 86.370 88.935 86.630 89.195 ;
        RECT 86.730 88.935 86.990 89.195 ;
        RECT 87.090 88.935 87.350 89.195 ;
        RECT 87.450 88.935 87.710 89.195 ;
        RECT 87.810 88.935 88.070 89.195 ;
        RECT 88.170 88.935 88.430 89.195 ;
        RECT 88.530 88.935 88.790 89.195 ;
        RECT 88.890 88.935 89.150 89.195 ;
        RECT 89.250 88.935 89.510 89.195 ;
        RECT 89.610 88.935 89.870 89.195 ;
        RECT 89.970 88.935 90.230 89.195 ;
        RECT 90.330 88.935 90.590 89.195 ;
        RECT 90.690 88.935 90.950 89.195 ;
        RECT 91.050 88.935 91.310 89.195 ;
        RECT 91.410 88.935 91.670 89.195 ;
        RECT 91.770 88.935 92.030 89.195 ;
        RECT 92.130 88.935 92.390 89.195 ;
        RECT 92.490 88.935 92.750 89.195 ;
        RECT 92.850 88.935 93.110 89.195 ;
        RECT 93.210 88.935 93.470 89.195 ;
        RECT 93.570 88.935 93.830 89.195 ;
        RECT 93.930 88.935 94.190 89.195 ;
        RECT 94.290 88.935 94.550 89.195 ;
        RECT 94.650 88.935 94.910 89.195 ;
        RECT 95.010 88.935 95.270 89.195 ;
        RECT 95.370 88.935 95.630 89.195 ;
        RECT 95.730 88.935 95.990 89.195 ;
        RECT 96.090 88.935 96.350 89.195 ;
        RECT 96.450 88.935 96.710 89.195 ;
        RECT 99.225 88.930 99.485 89.190 ;
        RECT 99.585 88.930 99.845 89.190 ;
        RECT 99.945 88.930 100.205 89.190 ;
        RECT 99.225 88.570 99.485 88.830 ;
        RECT 99.585 88.570 99.845 88.830 ;
        RECT 99.945 88.570 100.205 88.830 ;
        RECT 99.225 88.210 99.485 88.470 ;
        RECT 99.585 88.210 99.845 88.470 ;
        RECT 99.945 88.210 100.205 88.470 ;
        RECT 16.550 87.600 16.810 87.860 ;
        RECT 16.910 87.600 17.170 87.860 ;
        RECT 17.270 87.600 17.530 87.860 ;
        RECT 16.550 87.240 16.810 87.500 ;
        RECT 16.910 87.240 17.170 87.500 ;
        RECT 17.270 87.240 17.530 87.500 ;
        RECT 16.550 86.880 16.810 87.140 ;
        RECT 16.910 86.880 17.170 87.140 ;
        RECT 17.270 86.880 17.530 87.140 ;
        RECT 16.550 86.520 16.810 86.780 ;
        RECT 16.910 86.520 17.170 86.780 ;
        RECT 17.270 86.520 17.530 86.780 ;
        RECT 16.550 86.160 16.810 86.420 ;
        RECT 16.910 86.160 17.170 86.420 ;
        RECT 17.270 86.160 17.530 86.420 ;
        RECT 16.550 85.800 16.810 86.060 ;
        RECT 16.910 85.800 17.170 86.060 ;
        RECT 17.270 85.800 17.530 86.060 ;
        RECT 16.550 85.440 16.810 85.700 ;
        RECT 16.910 85.440 17.170 85.700 ;
        RECT 17.270 85.440 17.530 85.700 ;
        RECT 16.550 85.080 16.810 85.340 ;
        RECT 16.910 85.080 17.170 85.340 ;
        RECT 17.270 85.080 17.530 85.340 ;
        RECT 16.550 84.720 16.810 84.980 ;
        RECT 16.910 84.720 17.170 84.980 ;
        RECT 17.270 84.720 17.530 84.980 ;
        RECT 16.550 84.360 16.810 84.620 ;
        RECT 16.910 84.360 17.170 84.620 ;
        RECT 17.270 84.360 17.530 84.620 ;
        RECT 16.550 84.000 16.810 84.260 ;
        RECT 16.910 84.000 17.170 84.260 ;
        RECT 17.270 84.000 17.530 84.260 ;
        RECT 16.550 83.640 16.810 83.900 ;
        RECT 16.910 83.640 17.170 83.900 ;
        RECT 17.270 83.640 17.530 83.900 ;
        RECT 16.550 83.280 16.810 83.540 ;
        RECT 16.910 83.280 17.170 83.540 ;
        RECT 17.270 83.280 17.530 83.540 ;
        RECT 16.550 82.920 16.810 83.180 ;
        RECT 16.910 82.920 17.170 83.180 ;
        RECT 17.270 82.920 17.530 83.180 ;
        RECT 16.550 82.560 16.810 82.820 ;
        RECT 16.910 82.560 17.170 82.820 ;
        RECT 17.270 82.560 17.530 82.820 ;
        RECT 16.550 82.200 16.810 82.460 ;
        RECT 16.910 82.200 17.170 82.460 ;
        RECT 17.270 82.200 17.530 82.460 ;
        RECT 16.550 81.840 16.810 82.100 ;
        RECT 16.910 81.840 17.170 82.100 ;
        RECT 17.270 81.840 17.530 82.100 ;
        RECT 16.550 81.480 16.810 81.740 ;
        RECT 16.910 81.480 17.170 81.740 ;
        RECT 17.270 81.480 17.530 81.740 ;
        RECT 16.550 81.120 16.810 81.380 ;
        RECT 16.910 81.120 17.170 81.380 ;
        RECT 17.270 81.120 17.530 81.380 ;
        RECT 16.550 80.760 16.810 81.020 ;
        RECT 16.910 80.760 17.170 81.020 ;
        RECT 17.270 80.760 17.530 81.020 ;
        RECT 16.550 80.400 16.810 80.660 ;
        RECT 16.910 80.400 17.170 80.660 ;
        RECT 17.270 80.400 17.530 80.660 ;
        RECT 16.550 80.040 16.810 80.300 ;
        RECT 16.910 80.040 17.170 80.300 ;
        RECT 17.270 80.040 17.530 80.300 ;
        RECT 16.550 79.680 16.810 79.940 ;
        RECT 16.910 79.680 17.170 79.940 ;
        RECT 17.270 79.680 17.530 79.940 ;
        RECT 16.550 79.320 16.810 79.580 ;
        RECT 16.910 79.320 17.170 79.580 ;
        RECT 17.270 79.320 17.530 79.580 ;
        RECT 16.550 78.960 16.810 79.220 ;
        RECT 16.910 78.960 17.170 79.220 ;
        RECT 17.270 78.960 17.530 79.220 ;
        RECT 16.550 78.600 16.810 78.860 ;
        RECT 16.910 78.600 17.170 78.860 ;
        RECT 17.270 78.600 17.530 78.860 ;
        RECT 16.550 78.240 16.810 78.500 ;
        RECT 16.910 78.240 17.170 78.500 ;
        RECT 17.270 78.240 17.530 78.500 ;
        RECT 16.550 77.880 16.810 78.140 ;
        RECT 16.910 77.880 17.170 78.140 ;
        RECT 17.270 77.880 17.530 78.140 ;
        RECT 16.550 77.520 16.810 77.780 ;
        RECT 16.910 77.520 17.170 77.780 ;
        RECT 17.270 77.520 17.530 77.780 ;
        RECT 16.550 77.160 16.810 77.420 ;
        RECT 16.910 77.160 17.170 77.420 ;
        RECT 17.270 77.160 17.530 77.420 ;
        RECT 16.550 76.800 16.810 77.060 ;
        RECT 16.910 76.800 17.170 77.060 ;
        RECT 17.270 76.800 17.530 77.060 ;
        RECT 16.550 76.440 16.810 76.700 ;
        RECT 16.910 76.440 17.170 76.700 ;
        RECT 17.270 76.440 17.530 76.700 ;
        RECT 16.550 76.080 16.810 76.340 ;
        RECT 16.910 76.080 17.170 76.340 ;
        RECT 17.270 76.080 17.530 76.340 ;
        RECT 16.550 75.720 16.810 75.980 ;
        RECT 16.910 75.720 17.170 75.980 ;
        RECT 17.270 75.720 17.530 75.980 ;
        RECT 16.550 75.360 16.810 75.620 ;
        RECT 16.910 75.360 17.170 75.620 ;
        RECT 17.270 75.360 17.530 75.620 ;
        RECT 16.550 75.000 16.810 75.260 ;
        RECT 16.910 75.000 17.170 75.260 ;
        RECT 17.270 75.000 17.530 75.260 ;
        RECT 16.550 74.640 16.810 74.900 ;
        RECT 16.910 74.640 17.170 74.900 ;
        RECT 17.270 74.640 17.530 74.900 ;
        RECT 16.550 74.280 16.810 74.540 ;
        RECT 16.910 74.280 17.170 74.540 ;
        RECT 17.270 74.280 17.530 74.540 ;
        RECT 16.550 73.920 16.810 74.180 ;
        RECT 16.910 73.920 17.170 74.180 ;
        RECT 17.270 73.920 17.530 74.180 ;
        RECT 16.550 73.560 16.810 73.820 ;
        RECT 16.910 73.560 17.170 73.820 ;
        RECT 17.270 73.560 17.530 73.820 ;
        RECT 16.550 73.200 16.810 73.460 ;
        RECT 16.910 73.200 17.170 73.460 ;
        RECT 17.270 73.200 17.530 73.460 ;
        RECT 16.550 72.840 16.810 73.100 ;
        RECT 16.910 72.840 17.170 73.100 ;
        RECT 17.270 72.840 17.530 73.100 ;
        RECT 16.550 72.480 16.810 72.740 ;
        RECT 16.910 72.480 17.170 72.740 ;
        RECT 17.270 72.480 17.530 72.740 ;
        RECT 16.550 72.120 16.810 72.380 ;
        RECT 16.910 72.120 17.170 72.380 ;
        RECT 17.270 72.120 17.530 72.380 ;
        RECT 16.550 71.760 16.810 72.020 ;
        RECT 16.910 71.760 17.170 72.020 ;
        RECT 17.270 71.760 17.530 72.020 ;
        RECT 16.550 71.400 16.810 71.660 ;
        RECT 16.910 71.400 17.170 71.660 ;
        RECT 17.270 71.400 17.530 71.660 ;
        RECT 16.550 71.040 16.810 71.300 ;
        RECT 16.910 71.040 17.170 71.300 ;
        RECT 17.270 71.040 17.530 71.300 ;
        RECT 16.550 70.680 16.810 70.940 ;
        RECT 16.910 70.680 17.170 70.940 ;
        RECT 17.270 70.680 17.530 70.940 ;
        RECT 16.550 70.320 16.810 70.580 ;
        RECT 16.910 70.320 17.170 70.580 ;
        RECT 17.270 70.320 17.530 70.580 ;
        RECT 16.550 69.960 16.810 70.220 ;
        RECT 16.910 69.960 17.170 70.220 ;
        RECT 17.270 69.960 17.530 70.220 ;
        RECT 16.550 69.600 16.810 69.860 ;
        RECT 16.910 69.600 17.170 69.860 ;
        RECT 17.270 69.600 17.530 69.860 ;
        RECT 16.550 69.240 16.810 69.500 ;
        RECT 16.910 69.240 17.170 69.500 ;
        RECT 17.270 69.240 17.530 69.500 ;
        RECT 16.550 68.880 16.810 69.140 ;
        RECT 16.910 68.880 17.170 69.140 ;
        RECT 17.270 68.880 17.530 69.140 ;
        RECT 16.550 68.520 16.810 68.780 ;
        RECT 16.910 68.520 17.170 68.780 ;
        RECT 17.270 68.520 17.530 68.780 ;
        RECT 16.550 68.160 16.810 68.420 ;
        RECT 16.910 68.160 17.170 68.420 ;
        RECT 17.270 68.160 17.530 68.420 ;
        RECT 16.550 67.800 16.810 68.060 ;
        RECT 16.910 67.800 17.170 68.060 ;
        RECT 17.270 67.800 17.530 68.060 ;
        RECT 16.550 67.440 16.810 67.700 ;
        RECT 16.910 67.440 17.170 67.700 ;
        RECT 17.270 67.440 17.530 67.700 ;
        RECT 16.550 67.080 16.810 67.340 ;
        RECT 16.910 67.080 17.170 67.340 ;
        RECT 17.270 67.080 17.530 67.340 ;
        RECT 16.550 66.720 16.810 66.980 ;
        RECT 16.910 66.720 17.170 66.980 ;
        RECT 17.270 66.720 17.530 66.980 ;
        RECT 16.550 66.360 16.810 66.620 ;
        RECT 16.910 66.360 17.170 66.620 ;
        RECT 17.270 66.360 17.530 66.620 ;
        RECT 16.550 66.000 16.810 66.260 ;
        RECT 16.910 66.000 17.170 66.260 ;
        RECT 17.270 66.000 17.530 66.260 ;
        RECT 16.550 65.640 16.810 65.900 ;
        RECT 16.910 65.640 17.170 65.900 ;
        RECT 17.270 65.640 17.530 65.900 ;
        RECT 16.550 65.280 16.810 65.540 ;
        RECT 16.910 65.280 17.170 65.540 ;
        RECT 17.270 65.280 17.530 65.540 ;
        RECT 16.550 64.920 16.810 65.180 ;
        RECT 16.910 64.920 17.170 65.180 ;
        RECT 17.270 64.920 17.530 65.180 ;
        RECT 16.550 64.560 16.810 64.820 ;
        RECT 16.910 64.560 17.170 64.820 ;
        RECT 17.270 64.560 17.530 64.820 ;
        RECT 16.550 64.200 16.810 64.460 ;
        RECT 16.910 64.200 17.170 64.460 ;
        RECT 17.270 64.200 17.530 64.460 ;
        RECT 16.550 63.840 16.810 64.100 ;
        RECT 16.910 63.840 17.170 64.100 ;
        RECT 17.270 63.840 17.530 64.100 ;
        RECT 16.550 63.480 16.810 63.740 ;
        RECT 16.910 63.480 17.170 63.740 ;
        RECT 17.270 63.480 17.530 63.740 ;
        RECT 16.550 63.120 16.810 63.380 ;
        RECT 16.910 63.120 17.170 63.380 ;
        RECT 17.270 63.120 17.530 63.380 ;
        RECT 16.550 62.760 16.810 63.020 ;
        RECT 16.910 62.760 17.170 63.020 ;
        RECT 17.270 62.760 17.530 63.020 ;
        RECT 16.550 62.400 16.810 62.660 ;
        RECT 16.910 62.400 17.170 62.660 ;
        RECT 17.270 62.400 17.530 62.660 ;
        RECT 16.550 62.040 16.810 62.300 ;
        RECT 16.910 62.040 17.170 62.300 ;
        RECT 17.270 62.040 17.530 62.300 ;
        RECT 16.550 61.680 16.810 61.940 ;
        RECT 16.910 61.680 17.170 61.940 ;
        RECT 17.270 61.680 17.530 61.940 ;
        RECT 16.550 61.320 16.810 61.580 ;
        RECT 16.910 61.320 17.170 61.580 ;
        RECT 17.270 61.320 17.530 61.580 ;
        RECT 16.550 60.960 16.810 61.220 ;
        RECT 16.910 60.960 17.170 61.220 ;
        RECT 17.270 60.960 17.530 61.220 ;
        RECT 16.550 60.600 16.810 60.860 ;
        RECT 16.910 60.600 17.170 60.860 ;
        RECT 17.270 60.600 17.530 60.860 ;
        RECT 16.550 60.240 16.810 60.500 ;
        RECT 16.910 60.240 17.170 60.500 ;
        RECT 17.270 60.240 17.530 60.500 ;
        RECT 16.550 59.880 16.810 60.140 ;
        RECT 16.910 59.880 17.170 60.140 ;
        RECT 17.270 59.880 17.530 60.140 ;
        RECT 16.550 59.520 16.810 59.780 ;
        RECT 16.910 59.520 17.170 59.780 ;
        RECT 17.270 59.520 17.530 59.780 ;
        RECT 16.550 59.160 16.810 59.420 ;
        RECT 16.910 59.160 17.170 59.420 ;
        RECT 17.270 59.160 17.530 59.420 ;
        RECT 16.550 58.800 16.810 59.060 ;
        RECT 16.910 58.800 17.170 59.060 ;
        RECT 17.270 58.800 17.530 59.060 ;
        RECT 16.550 58.440 16.810 58.700 ;
        RECT 16.910 58.440 17.170 58.700 ;
        RECT 17.270 58.440 17.530 58.700 ;
        RECT 16.550 58.080 16.810 58.340 ;
        RECT 16.910 58.080 17.170 58.340 ;
        RECT 17.270 58.080 17.530 58.340 ;
        RECT 16.550 57.720 16.810 57.980 ;
        RECT 16.910 57.720 17.170 57.980 ;
        RECT 17.270 57.720 17.530 57.980 ;
        RECT 16.550 57.360 16.810 57.620 ;
        RECT 16.910 57.360 17.170 57.620 ;
        RECT 17.270 57.360 17.530 57.620 ;
        RECT 16.550 57.000 16.810 57.260 ;
        RECT 16.910 57.000 17.170 57.260 ;
        RECT 17.270 57.000 17.530 57.260 ;
        RECT 16.550 56.640 16.810 56.900 ;
        RECT 16.910 56.640 17.170 56.900 ;
        RECT 17.270 56.640 17.530 56.900 ;
        RECT 16.550 56.280 16.810 56.540 ;
        RECT 16.910 56.280 17.170 56.540 ;
        RECT 17.270 56.280 17.530 56.540 ;
        RECT 16.550 55.920 16.810 56.180 ;
        RECT 16.910 55.920 17.170 56.180 ;
        RECT 17.270 55.920 17.530 56.180 ;
        RECT 16.550 55.560 16.810 55.820 ;
        RECT 16.910 55.560 17.170 55.820 ;
        RECT 17.270 55.560 17.530 55.820 ;
        RECT 16.550 55.200 16.810 55.460 ;
        RECT 16.910 55.200 17.170 55.460 ;
        RECT 17.270 55.200 17.530 55.460 ;
        RECT 16.550 54.840 16.810 55.100 ;
        RECT 16.910 54.840 17.170 55.100 ;
        RECT 17.270 54.840 17.530 55.100 ;
        RECT 16.550 54.480 16.810 54.740 ;
        RECT 16.910 54.480 17.170 54.740 ;
        RECT 17.270 54.480 17.530 54.740 ;
        RECT 16.550 54.120 16.810 54.380 ;
        RECT 16.910 54.120 17.170 54.380 ;
        RECT 17.270 54.120 17.530 54.380 ;
        RECT 16.550 53.760 16.810 54.020 ;
        RECT 16.910 53.760 17.170 54.020 ;
        RECT 17.270 53.760 17.530 54.020 ;
        RECT 16.550 53.400 16.810 53.660 ;
        RECT 16.910 53.400 17.170 53.660 ;
        RECT 17.270 53.400 17.530 53.660 ;
        RECT 16.550 53.040 16.810 53.300 ;
        RECT 16.910 53.040 17.170 53.300 ;
        RECT 17.270 53.040 17.530 53.300 ;
        RECT 16.550 52.680 16.810 52.940 ;
        RECT 16.910 52.680 17.170 52.940 ;
        RECT 17.270 52.680 17.530 52.940 ;
        RECT 16.550 52.320 16.810 52.580 ;
        RECT 16.910 52.320 17.170 52.580 ;
        RECT 17.270 52.320 17.530 52.580 ;
        RECT 16.550 51.960 16.810 52.220 ;
        RECT 16.910 51.960 17.170 52.220 ;
        RECT 17.270 51.960 17.530 52.220 ;
        RECT 16.550 51.600 16.810 51.860 ;
        RECT 16.910 51.600 17.170 51.860 ;
        RECT 17.270 51.600 17.530 51.860 ;
        RECT 16.550 51.240 16.810 51.500 ;
        RECT 16.910 51.240 17.170 51.500 ;
        RECT 17.270 51.240 17.530 51.500 ;
        RECT 16.550 50.880 16.810 51.140 ;
        RECT 16.910 50.880 17.170 51.140 ;
        RECT 17.270 50.880 17.530 51.140 ;
        RECT 16.550 50.520 16.810 50.780 ;
        RECT 16.910 50.520 17.170 50.780 ;
        RECT 17.270 50.520 17.530 50.780 ;
        RECT 16.550 50.160 16.810 50.420 ;
        RECT 16.910 50.160 17.170 50.420 ;
        RECT 17.270 50.160 17.530 50.420 ;
        RECT 16.550 49.800 16.810 50.060 ;
        RECT 16.910 49.800 17.170 50.060 ;
        RECT 17.270 49.800 17.530 50.060 ;
        RECT 16.550 49.440 16.810 49.700 ;
        RECT 16.910 49.440 17.170 49.700 ;
        RECT 17.270 49.440 17.530 49.700 ;
        RECT 16.550 49.080 16.810 49.340 ;
        RECT 16.910 49.080 17.170 49.340 ;
        RECT 17.270 49.080 17.530 49.340 ;
        RECT 99.225 87.850 99.485 88.110 ;
        RECT 99.585 87.850 99.845 88.110 ;
        RECT 99.945 87.850 100.205 88.110 ;
        RECT 99.225 87.490 99.485 87.750 ;
        RECT 99.585 87.490 99.845 87.750 ;
        RECT 99.945 87.490 100.205 87.750 ;
        RECT 99.225 87.130 99.485 87.390 ;
        RECT 99.585 87.130 99.845 87.390 ;
        RECT 99.945 87.130 100.205 87.390 ;
        RECT 99.225 86.770 99.485 87.030 ;
        RECT 99.585 86.770 99.845 87.030 ;
        RECT 99.945 86.770 100.205 87.030 ;
        RECT 99.225 86.410 99.485 86.670 ;
        RECT 99.585 86.410 99.845 86.670 ;
        RECT 99.945 86.410 100.205 86.670 ;
        RECT 99.225 86.050 99.485 86.310 ;
        RECT 99.585 86.050 99.845 86.310 ;
        RECT 99.945 86.050 100.205 86.310 ;
        RECT 99.225 85.690 99.485 85.950 ;
        RECT 99.585 85.690 99.845 85.950 ;
        RECT 99.945 85.690 100.205 85.950 ;
        RECT 99.225 85.330 99.485 85.590 ;
        RECT 99.585 85.330 99.845 85.590 ;
        RECT 99.945 85.330 100.205 85.590 ;
        RECT 99.225 84.970 99.485 85.230 ;
        RECT 99.585 84.970 99.845 85.230 ;
        RECT 99.945 84.970 100.205 85.230 ;
        RECT 99.225 84.610 99.485 84.870 ;
        RECT 99.585 84.610 99.845 84.870 ;
        RECT 99.945 84.610 100.205 84.870 ;
        RECT 99.225 84.250 99.485 84.510 ;
        RECT 99.585 84.250 99.845 84.510 ;
        RECT 99.945 84.250 100.205 84.510 ;
        RECT 99.225 83.890 99.485 84.150 ;
        RECT 99.585 83.890 99.845 84.150 ;
        RECT 99.945 83.890 100.205 84.150 ;
        RECT 99.225 83.530 99.485 83.790 ;
        RECT 99.585 83.530 99.845 83.790 ;
        RECT 99.945 83.530 100.205 83.790 ;
        RECT 99.225 83.170 99.485 83.430 ;
        RECT 99.585 83.170 99.845 83.430 ;
        RECT 99.945 83.170 100.205 83.430 ;
        RECT 99.225 82.810 99.485 83.070 ;
        RECT 99.585 82.810 99.845 83.070 ;
        RECT 99.945 82.810 100.205 83.070 ;
        RECT 99.225 82.450 99.485 82.710 ;
        RECT 99.585 82.450 99.845 82.710 ;
        RECT 99.945 82.450 100.205 82.710 ;
        RECT 99.225 82.090 99.485 82.350 ;
        RECT 99.585 82.090 99.845 82.350 ;
        RECT 99.945 82.090 100.205 82.350 ;
        RECT 99.225 81.730 99.485 81.990 ;
        RECT 99.585 81.730 99.845 81.990 ;
        RECT 99.945 81.730 100.205 81.990 ;
        RECT 99.225 81.370 99.485 81.630 ;
        RECT 99.585 81.370 99.845 81.630 ;
        RECT 99.945 81.370 100.205 81.630 ;
        RECT 99.225 81.010 99.485 81.270 ;
        RECT 99.585 81.010 99.845 81.270 ;
        RECT 99.945 81.010 100.205 81.270 ;
        RECT 99.225 80.650 99.485 80.910 ;
        RECT 99.585 80.650 99.845 80.910 ;
        RECT 99.945 80.650 100.205 80.910 ;
        RECT 99.225 80.290 99.485 80.550 ;
        RECT 99.585 80.290 99.845 80.550 ;
        RECT 99.945 80.290 100.205 80.550 ;
        RECT 99.225 79.930 99.485 80.190 ;
        RECT 99.585 79.930 99.845 80.190 ;
        RECT 99.945 79.930 100.205 80.190 ;
        RECT 99.225 79.570 99.485 79.830 ;
        RECT 99.585 79.570 99.845 79.830 ;
        RECT 99.945 79.570 100.205 79.830 ;
        RECT 99.225 79.210 99.485 79.470 ;
        RECT 99.585 79.210 99.845 79.470 ;
        RECT 99.945 79.210 100.205 79.470 ;
        RECT 99.225 78.850 99.485 79.110 ;
        RECT 99.585 78.850 99.845 79.110 ;
        RECT 99.945 78.850 100.205 79.110 ;
        RECT 99.225 78.490 99.485 78.750 ;
        RECT 99.585 78.490 99.845 78.750 ;
        RECT 99.945 78.490 100.205 78.750 ;
        RECT 99.225 78.130 99.485 78.390 ;
        RECT 99.585 78.130 99.845 78.390 ;
        RECT 99.945 78.130 100.205 78.390 ;
        RECT 99.225 77.770 99.485 78.030 ;
        RECT 99.585 77.770 99.845 78.030 ;
        RECT 99.945 77.770 100.205 78.030 ;
        RECT 99.225 77.410 99.485 77.670 ;
        RECT 99.585 77.410 99.845 77.670 ;
        RECT 99.945 77.410 100.205 77.670 ;
        RECT 99.225 77.050 99.485 77.310 ;
        RECT 99.585 77.050 99.845 77.310 ;
        RECT 99.945 77.050 100.205 77.310 ;
        RECT 99.225 76.690 99.485 76.950 ;
        RECT 99.585 76.690 99.845 76.950 ;
        RECT 99.945 76.690 100.205 76.950 ;
        RECT 99.225 76.330 99.485 76.590 ;
        RECT 99.585 76.330 99.845 76.590 ;
        RECT 99.945 76.330 100.205 76.590 ;
        RECT 99.225 75.970 99.485 76.230 ;
        RECT 99.585 75.970 99.845 76.230 ;
        RECT 99.945 75.970 100.205 76.230 ;
        RECT 99.225 75.610 99.485 75.870 ;
        RECT 99.585 75.610 99.845 75.870 ;
        RECT 99.945 75.610 100.205 75.870 ;
        RECT 99.225 75.250 99.485 75.510 ;
        RECT 99.585 75.250 99.845 75.510 ;
        RECT 99.945 75.250 100.205 75.510 ;
        RECT 99.225 74.890 99.485 75.150 ;
        RECT 99.585 74.890 99.845 75.150 ;
        RECT 99.945 74.890 100.205 75.150 ;
        RECT 99.225 74.530 99.485 74.790 ;
        RECT 99.585 74.530 99.845 74.790 ;
        RECT 99.945 74.530 100.205 74.790 ;
        RECT 99.225 74.170 99.485 74.430 ;
        RECT 99.585 74.170 99.845 74.430 ;
        RECT 99.945 74.170 100.205 74.430 ;
        RECT 99.225 73.810 99.485 74.070 ;
        RECT 99.585 73.810 99.845 74.070 ;
        RECT 99.945 73.810 100.205 74.070 ;
        RECT 99.225 73.450 99.485 73.710 ;
        RECT 99.585 73.450 99.845 73.710 ;
        RECT 99.945 73.450 100.205 73.710 ;
        RECT 99.225 73.090 99.485 73.350 ;
        RECT 99.585 73.090 99.845 73.350 ;
        RECT 99.945 73.090 100.205 73.350 ;
        RECT 99.225 72.730 99.485 72.990 ;
        RECT 99.585 72.730 99.845 72.990 ;
        RECT 99.945 72.730 100.205 72.990 ;
        RECT 99.225 72.370 99.485 72.630 ;
        RECT 99.585 72.370 99.845 72.630 ;
        RECT 99.945 72.370 100.205 72.630 ;
        RECT 99.225 72.010 99.485 72.270 ;
        RECT 99.585 72.010 99.845 72.270 ;
        RECT 99.945 72.010 100.205 72.270 ;
        RECT 99.225 71.650 99.485 71.910 ;
        RECT 99.585 71.650 99.845 71.910 ;
        RECT 99.945 71.650 100.205 71.910 ;
        RECT 99.225 71.290 99.485 71.550 ;
        RECT 99.585 71.290 99.845 71.550 ;
        RECT 99.945 71.290 100.205 71.550 ;
        RECT 99.225 70.930 99.485 71.190 ;
        RECT 99.585 70.930 99.845 71.190 ;
        RECT 99.945 70.930 100.205 71.190 ;
        RECT 99.225 70.570 99.485 70.830 ;
        RECT 99.585 70.570 99.845 70.830 ;
        RECT 99.945 70.570 100.205 70.830 ;
        RECT 99.225 70.210 99.485 70.470 ;
        RECT 99.585 70.210 99.845 70.470 ;
        RECT 99.945 70.210 100.205 70.470 ;
        RECT 99.225 69.850 99.485 70.110 ;
        RECT 99.585 69.850 99.845 70.110 ;
        RECT 99.945 69.850 100.205 70.110 ;
        RECT 99.225 69.490 99.485 69.750 ;
        RECT 99.585 69.490 99.845 69.750 ;
        RECT 99.945 69.490 100.205 69.750 ;
        RECT 99.225 69.130 99.485 69.390 ;
        RECT 99.585 69.130 99.845 69.390 ;
        RECT 99.945 69.130 100.205 69.390 ;
        RECT 99.225 68.770 99.485 69.030 ;
        RECT 99.585 68.770 99.845 69.030 ;
        RECT 99.945 68.770 100.205 69.030 ;
        RECT 99.225 68.410 99.485 68.670 ;
        RECT 99.585 68.410 99.845 68.670 ;
        RECT 99.945 68.410 100.205 68.670 ;
        RECT 99.225 68.050 99.485 68.310 ;
        RECT 99.585 68.050 99.845 68.310 ;
        RECT 99.945 68.050 100.205 68.310 ;
        RECT 99.225 67.690 99.485 67.950 ;
        RECT 99.585 67.690 99.845 67.950 ;
        RECT 99.945 67.690 100.205 67.950 ;
        RECT 99.225 67.330 99.485 67.590 ;
        RECT 99.585 67.330 99.845 67.590 ;
        RECT 99.945 67.330 100.205 67.590 ;
        RECT 99.225 66.970 99.485 67.230 ;
        RECT 99.585 66.970 99.845 67.230 ;
        RECT 99.945 66.970 100.205 67.230 ;
        RECT 99.225 66.610 99.485 66.870 ;
        RECT 99.585 66.610 99.845 66.870 ;
        RECT 99.945 66.610 100.205 66.870 ;
        RECT 99.225 66.250 99.485 66.510 ;
        RECT 99.585 66.250 99.845 66.510 ;
        RECT 99.945 66.250 100.205 66.510 ;
        RECT 99.225 65.890 99.485 66.150 ;
        RECT 99.585 65.890 99.845 66.150 ;
        RECT 99.945 65.890 100.205 66.150 ;
        RECT 99.225 65.530 99.485 65.790 ;
        RECT 99.585 65.530 99.845 65.790 ;
        RECT 99.945 65.530 100.205 65.790 ;
        RECT 99.225 65.170 99.485 65.430 ;
        RECT 99.585 65.170 99.845 65.430 ;
        RECT 99.945 65.170 100.205 65.430 ;
        RECT 99.225 64.810 99.485 65.070 ;
        RECT 99.585 64.810 99.845 65.070 ;
        RECT 99.945 64.810 100.205 65.070 ;
        RECT 99.225 64.450 99.485 64.710 ;
        RECT 99.585 64.450 99.845 64.710 ;
        RECT 99.945 64.450 100.205 64.710 ;
        RECT 99.225 64.090 99.485 64.350 ;
        RECT 99.585 64.090 99.845 64.350 ;
        RECT 99.945 64.090 100.205 64.350 ;
        RECT 99.225 63.730 99.485 63.990 ;
        RECT 99.585 63.730 99.845 63.990 ;
        RECT 99.945 63.730 100.205 63.990 ;
        RECT 99.225 63.370 99.485 63.630 ;
        RECT 99.585 63.370 99.845 63.630 ;
        RECT 99.945 63.370 100.205 63.630 ;
        RECT 99.225 63.010 99.485 63.270 ;
        RECT 99.585 63.010 99.845 63.270 ;
        RECT 99.945 63.010 100.205 63.270 ;
        RECT 99.225 62.650 99.485 62.910 ;
        RECT 99.585 62.650 99.845 62.910 ;
        RECT 99.945 62.650 100.205 62.910 ;
        RECT 99.225 62.290 99.485 62.550 ;
        RECT 99.585 62.290 99.845 62.550 ;
        RECT 99.945 62.290 100.205 62.550 ;
        RECT 99.225 61.930 99.485 62.190 ;
        RECT 99.585 61.930 99.845 62.190 ;
        RECT 99.945 61.930 100.205 62.190 ;
        RECT 99.225 61.570 99.485 61.830 ;
        RECT 99.585 61.570 99.845 61.830 ;
        RECT 99.945 61.570 100.205 61.830 ;
        RECT 99.225 61.210 99.485 61.470 ;
        RECT 99.585 61.210 99.845 61.470 ;
        RECT 99.945 61.210 100.205 61.470 ;
        RECT 99.225 60.850 99.485 61.110 ;
        RECT 99.585 60.850 99.845 61.110 ;
        RECT 99.945 60.850 100.205 61.110 ;
        RECT 99.225 60.490 99.485 60.750 ;
        RECT 99.585 60.490 99.845 60.750 ;
        RECT 99.945 60.490 100.205 60.750 ;
        RECT 99.225 60.130 99.485 60.390 ;
        RECT 99.585 60.130 99.845 60.390 ;
        RECT 99.945 60.130 100.205 60.390 ;
        RECT 99.225 59.770 99.485 60.030 ;
        RECT 99.585 59.770 99.845 60.030 ;
        RECT 99.945 59.770 100.205 60.030 ;
        RECT 99.225 59.410 99.485 59.670 ;
        RECT 99.585 59.410 99.845 59.670 ;
        RECT 99.945 59.410 100.205 59.670 ;
        RECT 99.225 59.050 99.485 59.310 ;
        RECT 99.585 59.050 99.845 59.310 ;
        RECT 99.945 59.050 100.205 59.310 ;
        RECT 99.225 58.690 99.485 58.950 ;
        RECT 99.585 58.690 99.845 58.950 ;
        RECT 99.945 58.690 100.205 58.950 ;
        RECT 99.225 58.330 99.485 58.590 ;
        RECT 99.585 58.330 99.845 58.590 ;
        RECT 99.945 58.330 100.205 58.590 ;
        RECT 99.225 57.970 99.485 58.230 ;
        RECT 99.585 57.970 99.845 58.230 ;
        RECT 99.945 57.970 100.205 58.230 ;
        RECT 99.225 57.610 99.485 57.870 ;
        RECT 99.585 57.610 99.845 57.870 ;
        RECT 99.945 57.610 100.205 57.870 ;
        RECT 99.225 57.250 99.485 57.510 ;
        RECT 99.585 57.250 99.845 57.510 ;
        RECT 99.945 57.250 100.205 57.510 ;
        RECT 99.225 56.890 99.485 57.150 ;
        RECT 99.585 56.890 99.845 57.150 ;
        RECT 99.945 56.890 100.205 57.150 ;
        RECT 99.225 56.530 99.485 56.790 ;
        RECT 99.585 56.530 99.845 56.790 ;
        RECT 99.945 56.530 100.205 56.790 ;
        RECT 99.225 56.170 99.485 56.430 ;
        RECT 99.585 56.170 99.845 56.430 ;
        RECT 99.945 56.170 100.205 56.430 ;
        RECT 99.225 55.810 99.485 56.070 ;
        RECT 99.585 55.810 99.845 56.070 ;
        RECT 99.945 55.810 100.205 56.070 ;
        RECT 99.225 55.450 99.485 55.710 ;
        RECT 99.585 55.450 99.845 55.710 ;
        RECT 99.945 55.450 100.205 55.710 ;
        RECT 99.225 55.090 99.485 55.350 ;
        RECT 99.585 55.090 99.845 55.350 ;
        RECT 99.945 55.090 100.205 55.350 ;
        RECT 99.225 54.730 99.485 54.990 ;
        RECT 99.585 54.730 99.845 54.990 ;
        RECT 99.945 54.730 100.205 54.990 ;
        RECT 99.225 54.370 99.485 54.630 ;
        RECT 99.585 54.370 99.845 54.630 ;
        RECT 99.945 54.370 100.205 54.630 ;
        RECT 99.225 54.010 99.485 54.270 ;
        RECT 99.585 54.010 99.845 54.270 ;
        RECT 99.945 54.010 100.205 54.270 ;
        RECT 99.225 53.650 99.485 53.910 ;
        RECT 99.585 53.650 99.845 53.910 ;
        RECT 99.945 53.650 100.205 53.910 ;
        RECT 99.225 53.290 99.485 53.550 ;
        RECT 99.585 53.290 99.845 53.550 ;
        RECT 99.945 53.290 100.205 53.550 ;
        RECT 99.225 52.930 99.485 53.190 ;
        RECT 99.585 52.930 99.845 53.190 ;
        RECT 99.945 52.930 100.205 53.190 ;
        RECT 99.225 52.570 99.485 52.830 ;
        RECT 99.585 52.570 99.845 52.830 ;
        RECT 99.945 52.570 100.205 52.830 ;
        RECT 99.225 52.210 99.485 52.470 ;
        RECT 99.585 52.210 99.845 52.470 ;
        RECT 99.945 52.210 100.205 52.470 ;
        RECT 99.225 51.850 99.485 52.110 ;
        RECT 99.585 51.850 99.845 52.110 ;
        RECT 99.945 51.850 100.205 52.110 ;
        RECT 99.225 51.490 99.485 51.750 ;
        RECT 99.585 51.490 99.845 51.750 ;
        RECT 99.945 51.490 100.205 51.750 ;
        RECT 99.225 51.130 99.485 51.390 ;
        RECT 99.585 51.130 99.845 51.390 ;
        RECT 99.945 51.130 100.205 51.390 ;
        RECT 99.225 50.770 99.485 51.030 ;
        RECT 99.585 50.770 99.845 51.030 ;
        RECT 99.945 50.770 100.205 51.030 ;
        RECT 99.225 50.410 99.485 50.670 ;
        RECT 99.585 50.410 99.845 50.670 ;
        RECT 99.945 50.410 100.205 50.670 ;
        RECT 99.225 50.050 99.485 50.310 ;
        RECT 99.585 50.050 99.845 50.310 ;
        RECT 99.945 50.050 100.205 50.310 ;
        RECT 99.225 49.690 99.485 49.950 ;
        RECT 99.585 49.690 99.845 49.950 ;
        RECT 99.945 49.690 100.205 49.950 ;
        RECT 99.225 49.330 99.485 49.590 ;
        RECT 99.585 49.330 99.845 49.590 ;
        RECT 99.945 49.330 100.205 49.590 ;
        RECT 16.550 48.720 16.810 48.980 ;
        RECT 16.910 48.720 17.170 48.980 ;
        RECT 17.270 48.720 17.530 48.980 ;
        RECT 16.550 48.360 16.810 48.620 ;
        RECT 16.910 48.360 17.170 48.620 ;
        RECT 17.270 48.360 17.530 48.620 ;
        RECT 16.550 48.000 16.810 48.260 ;
        RECT 16.910 48.000 17.170 48.260 ;
        RECT 17.270 48.000 17.530 48.260 ;
        RECT 22.600 46.500 22.860 46.760 ;
        RECT 22.960 46.500 23.220 46.760 ;
        RECT 23.320 46.500 23.580 46.760 ;
        RECT 22.600 46.140 22.860 46.400 ;
        RECT 22.960 46.140 23.220 46.400 ;
        RECT 23.320 46.140 23.580 46.400 ;
        RECT 22.600 45.780 22.860 46.040 ;
        RECT 22.960 45.780 23.220 46.040 ;
        RECT 23.320 45.780 23.580 46.040 ;
        RECT 22.600 45.420 22.860 45.680 ;
        RECT 22.960 45.420 23.220 45.680 ;
        RECT 23.320 45.420 23.580 45.680 ;
        RECT 22.600 45.060 22.860 45.320 ;
        RECT 22.960 45.060 23.220 45.320 ;
        RECT 23.320 45.060 23.580 45.320 ;
        RECT 22.600 44.700 22.860 44.960 ;
        RECT 22.960 44.700 23.220 44.960 ;
        RECT 23.320 44.700 23.580 44.960 ;
        RECT 22.600 44.340 22.860 44.600 ;
        RECT 22.960 44.340 23.220 44.600 ;
        RECT 23.320 44.340 23.580 44.600 ;
        RECT 22.600 43.980 22.860 44.240 ;
        RECT 22.960 43.980 23.220 44.240 ;
        RECT 23.320 43.980 23.580 44.240 ;
        RECT 22.600 43.620 22.860 43.880 ;
        RECT 22.960 43.620 23.220 43.880 ;
        RECT 23.320 43.620 23.580 43.880 ;
        RECT 22.600 43.260 22.860 43.520 ;
        RECT 22.960 43.260 23.220 43.520 ;
        RECT 23.320 43.260 23.580 43.520 ;
        RECT 22.600 42.900 22.860 43.160 ;
        RECT 22.960 42.900 23.220 43.160 ;
        RECT 23.320 42.900 23.580 43.160 ;
        RECT 22.600 42.540 22.860 42.800 ;
        RECT 22.960 42.540 23.220 42.800 ;
        RECT 23.320 42.540 23.580 42.800 ;
        RECT 22.600 42.180 22.860 42.440 ;
        RECT 22.960 42.180 23.220 42.440 ;
        RECT 23.320 42.180 23.580 42.440 ;
        RECT 22.600 41.820 22.860 42.080 ;
        RECT 22.960 41.820 23.220 42.080 ;
        RECT 23.320 41.820 23.580 42.080 ;
        RECT 22.600 41.460 22.860 41.720 ;
        RECT 22.960 41.460 23.220 41.720 ;
        RECT 23.320 41.460 23.580 41.720 ;
        RECT 22.600 41.100 22.860 41.360 ;
        RECT 22.960 41.100 23.220 41.360 ;
        RECT 23.320 41.100 23.580 41.360 ;
        RECT 22.600 40.740 22.860 41.000 ;
        RECT 22.960 40.740 23.220 41.000 ;
        RECT 23.320 40.740 23.580 41.000 ;
        RECT 22.600 40.380 22.860 40.640 ;
        RECT 22.960 40.380 23.220 40.640 ;
        RECT 23.320 40.380 23.580 40.640 ;
        RECT 22.600 40.020 22.860 40.280 ;
        RECT 22.960 40.020 23.220 40.280 ;
        RECT 23.320 40.020 23.580 40.280 ;
        RECT 22.600 39.660 22.860 39.920 ;
        RECT 22.960 39.660 23.220 39.920 ;
        RECT 23.320 39.660 23.580 39.920 ;
        RECT 22.600 39.300 22.860 39.560 ;
        RECT 22.960 39.300 23.220 39.560 ;
        RECT 23.320 39.300 23.580 39.560 ;
        RECT 22.600 38.940 22.860 39.200 ;
        RECT 22.960 38.940 23.220 39.200 ;
        RECT 23.320 38.940 23.580 39.200 ;
        RECT 22.600 38.580 22.860 38.840 ;
        RECT 22.960 38.580 23.220 38.840 ;
        RECT 23.320 38.580 23.580 38.840 ;
        RECT 22.600 38.220 22.860 38.480 ;
        RECT 22.960 38.220 23.220 38.480 ;
        RECT 23.320 38.220 23.580 38.480 ;
        RECT 22.600 37.860 22.860 38.120 ;
        RECT 22.960 37.860 23.220 38.120 ;
        RECT 23.320 37.860 23.580 38.120 ;
        RECT 22.600 37.500 22.860 37.760 ;
        RECT 22.960 37.500 23.220 37.760 ;
        RECT 23.320 37.500 23.580 37.760 ;
        RECT 22.600 37.140 22.860 37.400 ;
        RECT 22.960 37.140 23.220 37.400 ;
        RECT 23.320 37.140 23.580 37.400 ;
        RECT 22.600 36.780 22.860 37.040 ;
        RECT 22.960 36.780 23.220 37.040 ;
        RECT 23.320 36.780 23.580 37.040 ;
        RECT 22.600 36.420 22.860 36.680 ;
        RECT 22.960 36.420 23.220 36.680 ;
        RECT 23.320 36.420 23.580 36.680 ;
        RECT 22.600 36.060 22.860 36.320 ;
        RECT 22.960 36.060 23.220 36.320 ;
        RECT 23.320 36.060 23.580 36.320 ;
        RECT 22.600 35.700 22.860 35.960 ;
        RECT 22.960 35.700 23.220 35.960 ;
        RECT 23.320 35.700 23.580 35.960 ;
        RECT 22.600 35.340 22.860 35.600 ;
        RECT 22.960 35.340 23.220 35.600 ;
        RECT 23.320 35.340 23.580 35.600 ;
        RECT 22.600 34.980 22.860 35.240 ;
        RECT 22.960 34.980 23.220 35.240 ;
        RECT 23.320 34.980 23.580 35.240 ;
        RECT 22.600 34.620 22.860 34.880 ;
        RECT 22.960 34.620 23.220 34.880 ;
        RECT 23.320 34.620 23.580 34.880 ;
        RECT 22.600 34.260 22.860 34.520 ;
        RECT 22.960 34.260 23.220 34.520 ;
        RECT 23.320 34.260 23.580 34.520 ;
        RECT 22.600 33.900 22.860 34.160 ;
        RECT 22.960 33.900 23.220 34.160 ;
        RECT 23.320 33.900 23.580 34.160 ;
        RECT 22.600 33.540 22.860 33.800 ;
        RECT 22.960 33.540 23.220 33.800 ;
        RECT 23.320 33.540 23.580 33.800 ;
        RECT 22.600 33.180 22.860 33.440 ;
        RECT 22.960 33.180 23.220 33.440 ;
        RECT 23.320 33.180 23.580 33.440 ;
        RECT 22.600 32.820 22.860 33.080 ;
        RECT 22.960 32.820 23.220 33.080 ;
        RECT 23.320 32.820 23.580 33.080 ;
        RECT 22.600 32.460 22.860 32.720 ;
        RECT 22.960 32.460 23.220 32.720 ;
        RECT 23.320 32.460 23.580 32.720 ;
        RECT 22.600 32.100 22.860 32.360 ;
        RECT 22.960 32.100 23.220 32.360 ;
        RECT 23.320 32.100 23.580 32.360 ;
        RECT 22.600 31.740 22.860 32.000 ;
        RECT 22.960 31.740 23.220 32.000 ;
        RECT 23.320 31.740 23.580 32.000 ;
        RECT 22.600 31.380 22.860 31.640 ;
        RECT 22.960 31.380 23.220 31.640 ;
        RECT 23.320 31.380 23.580 31.640 ;
        RECT 22.600 31.020 22.860 31.280 ;
        RECT 22.960 31.020 23.220 31.280 ;
        RECT 23.320 31.020 23.580 31.280 ;
        RECT 22.600 30.660 22.860 30.920 ;
        RECT 22.960 30.660 23.220 30.920 ;
        RECT 23.320 30.660 23.580 30.920 ;
        RECT 22.600 30.300 22.860 30.560 ;
        RECT 22.960 30.300 23.220 30.560 ;
        RECT 23.320 30.300 23.580 30.560 ;
        RECT 22.600 29.940 22.860 30.200 ;
        RECT 22.960 29.940 23.220 30.200 ;
        RECT 23.320 29.940 23.580 30.200 ;
        RECT 22.600 29.580 22.860 29.840 ;
        RECT 22.960 29.580 23.220 29.840 ;
        RECT 23.320 29.580 23.580 29.840 ;
        RECT 22.600 29.220 22.860 29.480 ;
        RECT 22.960 29.220 23.220 29.480 ;
        RECT 23.320 29.220 23.580 29.480 ;
        RECT 22.600 28.860 22.860 29.120 ;
        RECT 22.960 28.860 23.220 29.120 ;
        RECT 23.320 28.860 23.580 29.120 ;
        RECT 22.600 28.500 22.860 28.760 ;
        RECT 22.960 28.500 23.220 28.760 ;
        RECT 23.320 28.500 23.580 28.760 ;
        RECT 22.600 28.140 22.860 28.400 ;
        RECT 22.960 28.140 23.220 28.400 ;
        RECT 23.320 28.140 23.580 28.400 ;
        RECT 22.600 27.780 22.860 28.040 ;
        RECT 22.960 27.780 23.220 28.040 ;
        RECT 23.320 27.780 23.580 28.040 ;
        RECT 22.600 27.420 22.860 27.680 ;
        RECT 22.960 27.420 23.220 27.680 ;
        RECT 23.320 27.420 23.580 27.680 ;
        RECT 22.600 27.060 22.860 27.320 ;
        RECT 22.960 27.060 23.220 27.320 ;
        RECT 23.320 27.060 23.580 27.320 ;
        RECT 22.600 26.700 22.860 26.960 ;
        RECT 22.960 26.700 23.220 26.960 ;
        RECT 23.320 26.700 23.580 26.960 ;
        RECT 65.255 27.605 65.515 27.865 ;
        RECT 65.615 27.605 65.875 27.865 ;
        RECT 65.975 27.605 66.235 27.865 ;
        RECT 66.335 27.605 66.595 27.865 ;
        RECT 66.695 27.605 66.955 27.865 ;
        RECT 67.055 27.605 67.315 27.865 ;
        RECT 67.415 27.605 67.675 27.865 ;
        RECT 67.775 27.605 68.035 27.865 ;
        RECT 68.135 27.605 68.395 27.865 ;
        RECT 68.495 27.605 68.755 27.865 ;
        RECT 68.855 27.605 69.115 27.865 ;
        RECT 69.215 27.605 69.475 27.865 ;
        RECT 69.575 27.605 69.835 27.865 ;
        RECT 69.935 27.605 70.195 27.865 ;
        RECT 70.295 27.605 70.555 27.865 ;
        RECT 70.655 27.605 70.915 27.865 ;
        RECT 71.015 27.605 71.275 27.865 ;
        RECT 71.375 27.605 71.635 27.865 ;
        RECT 71.735 27.605 71.995 27.865 ;
        RECT 72.095 27.605 72.355 27.865 ;
        RECT 72.455 27.605 72.715 27.865 ;
        RECT 72.815 27.605 73.075 27.865 ;
        RECT 73.175 27.605 73.435 27.865 ;
        RECT 73.535 27.605 73.795 27.865 ;
        RECT 73.895 27.605 74.155 27.865 ;
        RECT 74.255 27.605 74.515 27.865 ;
        RECT 74.615 27.605 74.875 27.865 ;
        RECT 74.975 27.605 75.235 27.865 ;
        RECT 75.335 27.605 75.595 27.865 ;
        RECT 75.695 27.605 75.955 27.865 ;
        RECT 76.055 27.605 76.315 27.865 ;
        RECT 76.415 27.605 76.675 27.865 ;
        RECT 76.775 27.605 77.035 27.865 ;
        RECT 77.135 27.605 77.395 27.865 ;
        RECT 77.495 27.605 77.755 27.865 ;
        RECT 77.855 27.605 78.115 27.865 ;
        RECT 78.215 27.605 78.475 27.865 ;
        RECT 78.575 27.605 78.835 27.865 ;
        RECT 78.935 27.605 79.195 27.865 ;
        RECT 79.295 27.605 79.555 27.865 ;
        RECT 79.655 27.605 79.915 27.865 ;
        RECT 80.015 27.605 80.275 27.865 ;
        RECT 80.375 27.605 80.635 27.865 ;
        RECT 80.735 27.605 80.995 27.865 ;
        RECT 81.095 27.605 81.355 27.865 ;
        RECT 81.455 27.605 81.715 27.865 ;
        RECT 81.815 27.605 82.075 27.865 ;
        RECT 82.175 27.605 82.435 27.865 ;
        RECT 82.535 27.605 82.795 27.865 ;
        RECT 82.895 27.605 83.155 27.865 ;
        RECT 83.255 27.605 83.515 27.865 ;
        RECT 83.615 27.605 83.875 27.865 ;
        RECT 83.975 27.605 84.235 27.865 ;
        RECT 84.335 27.605 84.595 27.865 ;
        RECT 84.695 27.605 84.955 27.865 ;
        RECT 85.055 27.605 85.315 27.865 ;
        RECT 85.415 27.605 85.675 27.865 ;
        RECT 85.775 27.605 86.035 27.865 ;
        RECT 86.135 27.605 86.395 27.865 ;
        RECT 86.495 27.605 86.755 27.865 ;
        RECT 86.855 27.605 87.115 27.865 ;
        RECT 87.215 27.605 87.475 27.865 ;
        RECT 87.575 27.605 87.835 27.865 ;
        RECT 87.935 27.605 88.195 27.865 ;
        RECT 88.295 27.605 88.555 27.865 ;
        RECT 88.655 27.605 88.915 27.865 ;
        RECT 89.015 27.605 89.275 27.865 ;
        RECT 89.375 27.605 89.635 27.865 ;
        RECT 89.735 27.605 89.995 27.865 ;
        RECT 90.095 27.605 90.355 27.865 ;
        RECT 90.455 27.605 90.715 27.865 ;
        RECT 90.815 27.605 91.075 27.865 ;
        RECT 91.175 27.605 91.435 27.865 ;
        RECT 91.535 27.605 91.795 27.865 ;
        RECT 91.895 27.605 92.155 27.865 ;
        RECT 92.255 27.605 92.515 27.865 ;
        RECT 92.615 27.605 92.875 27.865 ;
        RECT 92.975 27.605 93.235 27.865 ;
        RECT 93.335 27.605 93.595 27.865 ;
        RECT 93.695 27.605 93.955 27.865 ;
        RECT 94.055 27.605 94.315 27.865 ;
        RECT 94.415 27.605 94.675 27.865 ;
        RECT 94.775 27.605 95.035 27.865 ;
        RECT 95.135 27.605 95.395 27.865 ;
        RECT 95.495 27.605 95.755 27.865 ;
        RECT 95.855 27.605 96.115 27.865 ;
        RECT 96.215 27.605 96.475 27.865 ;
        RECT 96.575 27.605 96.835 27.865 ;
        RECT 96.935 27.605 97.195 27.865 ;
        RECT 97.295 27.605 97.555 27.865 ;
        RECT 97.655 27.605 97.915 27.865 ;
        RECT 98.015 27.605 98.275 27.865 ;
        RECT 98.375 27.605 98.635 27.865 ;
        RECT 98.735 27.605 98.995 27.865 ;
        RECT 99.095 27.605 99.355 27.865 ;
        RECT 99.455 27.605 99.715 27.865 ;
        RECT 99.815 27.605 100.075 27.865 ;
        RECT 100.175 27.605 100.435 27.865 ;
        RECT 100.535 27.605 100.795 27.865 ;
        RECT 100.895 27.605 101.155 27.865 ;
        RECT 101.255 27.605 101.515 27.865 ;
        RECT 101.615 27.605 101.875 27.865 ;
        RECT 101.975 27.605 102.235 27.865 ;
        RECT 102.335 27.605 102.595 27.865 ;
        RECT 102.695 27.605 102.955 27.865 ;
        RECT 103.055 27.605 103.315 27.865 ;
        RECT 103.415 27.605 103.675 27.865 ;
        RECT 103.775 27.605 104.035 27.865 ;
        RECT 104.135 27.605 104.395 27.865 ;
        RECT 104.495 27.605 104.755 27.865 ;
        RECT 104.855 27.605 105.115 27.865 ;
        RECT 65.255 27.245 65.515 27.505 ;
        RECT 65.615 27.245 65.875 27.505 ;
        RECT 65.975 27.245 66.235 27.505 ;
        RECT 66.335 27.245 66.595 27.505 ;
        RECT 66.695 27.245 66.955 27.505 ;
        RECT 67.055 27.245 67.315 27.505 ;
        RECT 67.415 27.245 67.675 27.505 ;
        RECT 67.775 27.245 68.035 27.505 ;
        RECT 68.135 27.245 68.395 27.505 ;
        RECT 68.495 27.245 68.755 27.505 ;
        RECT 68.855 27.245 69.115 27.505 ;
        RECT 69.215 27.245 69.475 27.505 ;
        RECT 69.575 27.245 69.835 27.505 ;
        RECT 69.935 27.245 70.195 27.505 ;
        RECT 70.295 27.245 70.555 27.505 ;
        RECT 70.655 27.245 70.915 27.505 ;
        RECT 71.015 27.245 71.275 27.505 ;
        RECT 71.375 27.245 71.635 27.505 ;
        RECT 71.735 27.245 71.995 27.505 ;
        RECT 72.095 27.245 72.355 27.505 ;
        RECT 72.455 27.245 72.715 27.505 ;
        RECT 72.815 27.245 73.075 27.505 ;
        RECT 73.175 27.245 73.435 27.505 ;
        RECT 73.535 27.245 73.795 27.505 ;
        RECT 73.895 27.245 74.155 27.505 ;
        RECT 74.255 27.245 74.515 27.505 ;
        RECT 74.615 27.245 74.875 27.505 ;
        RECT 74.975 27.245 75.235 27.505 ;
        RECT 75.335 27.245 75.595 27.505 ;
        RECT 75.695 27.245 75.955 27.505 ;
        RECT 76.055 27.245 76.315 27.505 ;
        RECT 76.415 27.245 76.675 27.505 ;
        RECT 76.775 27.245 77.035 27.505 ;
        RECT 77.135 27.245 77.395 27.505 ;
        RECT 77.495 27.245 77.755 27.505 ;
        RECT 77.855 27.245 78.115 27.505 ;
        RECT 78.215 27.245 78.475 27.505 ;
        RECT 78.575 27.245 78.835 27.505 ;
        RECT 78.935 27.245 79.195 27.505 ;
        RECT 79.295 27.245 79.555 27.505 ;
        RECT 79.655 27.245 79.915 27.505 ;
        RECT 80.015 27.245 80.275 27.505 ;
        RECT 80.375 27.245 80.635 27.505 ;
        RECT 80.735 27.245 80.995 27.505 ;
        RECT 81.095 27.245 81.355 27.505 ;
        RECT 81.455 27.245 81.715 27.505 ;
        RECT 81.815 27.245 82.075 27.505 ;
        RECT 82.175 27.245 82.435 27.505 ;
        RECT 82.535 27.245 82.795 27.505 ;
        RECT 82.895 27.245 83.155 27.505 ;
        RECT 83.255 27.245 83.515 27.505 ;
        RECT 83.615 27.245 83.875 27.505 ;
        RECT 83.975 27.245 84.235 27.505 ;
        RECT 84.335 27.245 84.595 27.505 ;
        RECT 84.695 27.245 84.955 27.505 ;
        RECT 85.055 27.245 85.315 27.505 ;
        RECT 85.415 27.245 85.675 27.505 ;
        RECT 85.775 27.245 86.035 27.505 ;
        RECT 86.135 27.245 86.395 27.505 ;
        RECT 86.495 27.245 86.755 27.505 ;
        RECT 86.855 27.245 87.115 27.505 ;
        RECT 87.215 27.245 87.475 27.505 ;
        RECT 87.575 27.245 87.835 27.505 ;
        RECT 87.935 27.245 88.195 27.505 ;
        RECT 88.295 27.245 88.555 27.505 ;
        RECT 88.655 27.245 88.915 27.505 ;
        RECT 89.015 27.245 89.275 27.505 ;
        RECT 89.375 27.245 89.635 27.505 ;
        RECT 89.735 27.245 89.995 27.505 ;
        RECT 90.095 27.245 90.355 27.505 ;
        RECT 90.455 27.245 90.715 27.505 ;
        RECT 90.815 27.245 91.075 27.505 ;
        RECT 91.175 27.245 91.435 27.505 ;
        RECT 91.535 27.245 91.795 27.505 ;
        RECT 91.895 27.245 92.155 27.505 ;
        RECT 92.255 27.245 92.515 27.505 ;
        RECT 92.615 27.245 92.875 27.505 ;
        RECT 92.975 27.245 93.235 27.505 ;
        RECT 93.335 27.245 93.595 27.505 ;
        RECT 93.695 27.245 93.955 27.505 ;
        RECT 94.055 27.245 94.315 27.505 ;
        RECT 94.415 27.245 94.675 27.505 ;
        RECT 94.775 27.245 95.035 27.505 ;
        RECT 95.135 27.245 95.395 27.505 ;
        RECT 95.495 27.245 95.755 27.505 ;
        RECT 95.855 27.245 96.115 27.505 ;
        RECT 96.215 27.245 96.475 27.505 ;
        RECT 96.575 27.245 96.835 27.505 ;
        RECT 96.935 27.245 97.195 27.505 ;
        RECT 97.295 27.245 97.555 27.505 ;
        RECT 97.655 27.245 97.915 27.505 ;
        RECT 98.015 27.245 98.275 27.505 ;
        RECT 98.375 27.245 98.635 27.505 ;
        RECT 98.735 27.245 98.995 27.505 ;
        RECT 99.095 27.245 99.355 27.505 ;
        RECT 99.455 27.245 99.715 27.505 ;
        RECT 99.815 27.245 100.075 27.505 ;
        RECT 100.175 27.245 100.435 27.505 ;
        RECT 100.535 27.245 100.795 27.505 ;
        RECT 100.895 27.245 101.155 27.505 ;
        RECT 101.255 27.245 101.515 27.505 ;
        RECT 101.615 27.245 101.875 27.505 ;
        RECT 101.975 27.245 102.235 27.505 ;
        RECT 102.335 27.245 102.595 27.505 ;
        RECT 102.695 27.245 102.955 27.505 ;
        RECT 103.055 27.245 103.315 27.505 ;
        RECT 103.415 27.245 103.675 27.505 ;
        RECT 103.775 27.245 104.035 27.505 ;
        RECT 104.135 27.245 104.395 27.505 ;
        RECT 104.495 27.245 104.755 27.505 ;
        RECT 104.855 27.245 105.115 27.505 ;
        RECT 22.600 26.340 22.860 26.600 ;
        RECT 22.960 26.340 23.220 26.600 ;
        RECT 23.320 26.340 23.580 26.600 ;
        RECT 22.600 25.980 22.860 26.240 ;
        RECT 22.960 25.980 23.220 26.240 ;
        RECT 23.320 25.980 23.580 26.240 ;
        RECT 22.600 25.620 22.860 25.880 ;
        RECT 22.960 25.620 23.220 25.880 ;
        RECT 23.320 25.620 23.580 25.880 ;
        RECT 65.255 26.885 65.515 27.145 ;
        RECT 65.615 26.885 65.875 27.145 ;
        RECT 65.975 26.885 66.235 27.145 ;
        RECT 66.335 26.885 66.595 27.145 ;
        RECT 66.695 26.885 66.955 27.145 ;
        RECT 67.055 26.885 67.315 27.145 ;
        RECT 67.415 26.885 67.675 27.145 ;
        RECT 67.775 26.885 68.035 27.145 ;
        RECT 68.135 26.885 68.395 27.145 ;
        RECT 68.495 26.885 68.755 27.145 ;
        RECT 68.855 26.885 69.115 27.145 ;
        RECT 69.215 26.885 69.475 27.145 ;
        RECT 69.575 26.885 69.835 27.145 ;
        RECT 69.935 26.885 70.195 27.145 ;
        RECT 70.295 26.885 70.555 27.145 ;
        RECT 70.655 26.885 70.915 27.145 ;
        RECT 71.015 26.885 71.275 27.145 ;
        RECT 71.375 26.885 71.635 27.145 ;
        RECT 71.735 26.885 71.995 27.145 ;
        RECT 72.095 26.885 72.355 27.145 ;
        RECT 72.455 26.885 72.715 27.145 ;
        RECT 72.815 26.885 73.075 27.145 ;
        RECT 73.175 26.885 73.435 27.145 ;
        RECT 73.535 26.885 73.795 27.145 ;
        RECT 73.895 26.885 74.155 27.145 ;
        RECT 74.255 26.885 74.515 27.145 ;
        RECT 74.615 26.885 74.875 27.145 ;
        RECT 74.975 26.885 75.235 27.145 ;
        RECT 75.335 26.885 75.595 27.145 ;
        RECT 75.695 26.885 75.955 27.145 ;
        RECT 76.055 26.885 76.315 27.145 ;
        RECT 76.415 26.885 76.675 27.145 ;
        RECT 76.775 26.885 77.035 27.145 ;
        RECT 77.135 26.885 77.395 27.145 ;
        RECT 77.495 26.885 77.755 27.145 ;
        RECT 77.855 26.885 78.115 27.145 ;
        RECT 78.215 26.885 78.475 27.145 ;
        RECT 78.575 26.885 78.835 27.145 ;
        RECT 78.935 26.885 79.195 27.145 ;
        RECT 79.295 26.885 79.555 27.145 ;
        RECT 79.655 26.885 79.915 27.145 ;
        RECT 80.015 26.885 80.275 27.145 ;
        RECT 80.375 26.885 80.635 27.145 ;
        RECT 80.735 26.885 80.995 27.145 ;
        RECT 81.095 26.885 81.355 27.145 ;
        RECT 81.455 26.885 81.715 27.145 ;
        RECT 81.815 26.885 82.075 27.145 ;
        RECT 82.175 26.885 82.435 27.145 ;
        RECT 82.535 26.885 82.795 27.145 ;
        RECT 82.895 26.885 83.155 27.145 ;
        RECT 83.255 26.885 83.515 27.145 ;
        RECT 83.615 26.885 83.875 27.145 ;
        RECT 83.975 26.885 84.235 27.145 ;
        RECT 84.335 26.885 84.595 27.145 ;
        RECT 84.695 26.885 84.955 27.145 ;
        RECT 85.055 26.885 85.315 27.145 ;
        RECT 85.415 26.885 85.675 27.145 ;
        RECT 85.775 26.885 86.035 27.145 ;
        RECT 86.135 26.885 86.395 27.145 ;
        RECT 86.495 26.885 86.755 27.145 ;
        RECT 86.855 26.885 87.115 27.145 ;
        RECT 87.215 26.885 87.475 27.145 ;
        RECT 87.575 26.885 87.835 27.145 ;
        RECT 87.935 26.885 88.195 27.145 ;
        RECT 88.295 26.885 88.555 27.145 ;
        RECT 88.655 26.885 88.915 27.145 ;
        RECT 89.015 26.885 89.275 27.145 ;
        RECT 89.375 26.885 89.635 27.145 ;
        RECT 89.735 26.885 89.995 27.145 ;
        RECT 90.095 26.885 90.355 27.145 ;
        RECT 90.455 26.885 90.715 27.145 ;
        RECT 90.815 26.885 91.075 27.145 ;
        RECT 91.175 26.885 91.435 27.145 ;
        RECT 91.535 26.885 91.795 27.145 ;
        RECT 91.895 26.885 92.155 27.145 ;
        RECT 92.255 26.885 92.515 27.145 ;
        RECT 92.615 26.885 92.875 27.145 ;
        RECT 92.975 26.885 93.235 27.145 ;
        RECT 93.335 26.885 93.595 27.145 ;
        RECT 93.695 26.885 93.955 27.145 ;
        RECT 94.055 26.885 94.315 27.145 ;
        RECT 94.415 26.885 94.675 27.145 ;
        RECT 94.775 26.885 95.035 27.145 ;
        RECT 95.135 26.885 95.395 27.145 ;
        RECT 95.495 26.885 95.755 27.145 ;
        RECT 95.855 26.885 96.115 27.145 ;
        RECT 96.215 26.885 96.475 27.145 ;
        RECT 96.575 26.885 96.835 27.145 ;
        RECT 96.935 26.885 97.195 27.145 ;
        RECT 97.295 26.885 97.555 27.145 ;
        RECT 97.655 26.885 97.915 27.145 ;
        RECT 98.015 26.885 98.275 27.145 ;
        RECT 98.375 26.885 98.635 27.145 ;
        RECT 98.735 26.885 98.995 27.145 ;
        RECT 99.095 26.885 99.355 27.145 ;
        RECT 99.455 26.885 99.715 27.145 ;
        RECT 99.815 26.885 100.075 27.145 ;
        RECT 100.175 26.885 100.435 27.145 ;
        RECT 100.535 26.885 100.795 27.145 ;
        RECT 100.895 26.885 101.155 27.145 ;
        RECT 101.255 26.885 101.515 27.145 ;
        RECT 101.615 26.885 101.875 27.145 ;
        RECT 101.975 26.885 102.235 27.145 ;
        RECT 102.335 26.885 102.595 27.145 ;
        RECT 102.695 26.885 102.955 27.145 ;
        RECT 103.055 26.885 103.315 27.145 ;
        RECT 103.415 26.885 103.675 27.145 ;
        RECT 103.775 26.885 104.035 27.145 ;
        RECT 104.135 26.885 104.395 27.145 ;
        RECT 104.495 26.885 104.755 27.145 ;
        RECT 104.855 26.885 105.115 27.145 ;
        RECT 22.600 25.260 22.860 25.520 ;
        RECT 22.960 25.260 23.220 25.520 ;
        RECT 23.320 25.260 23.580 25.520 ;
        RECT 22.600 24.900 22.860 25.160 ;
        RECT 22.960 24.900 23.220 25.160 ;
        RECT 23.320 24.900 23.580 25.160 ;
        RECT 22.600 24.540 22.860 24.800 ;
        RECT 22.960 24.540 23.220 24.800 ;
        RECT 23.320 24.540 23.580 24.800 ;
        RECT 22.600 24.180 22.860 24.440 ;
        RECT 22.960 24.180 23.220 24.440 ;
        RECT 23.320 24.180 23.580 24.440 ;
        RECT 22.600 23.820 22.860 24.080 ;
        RECT 22.960 23.820 23.220 24.080 ;
        RECT 23.320 23.820 23.580 24.080 ;
        RECT 22.600 23.460 22.860 23.720 ;
        RECT 22.960 23.460 23.220 23.720 ;
        RECT 23.320 23.460 23.580 23.720 ;
        RECT 22.600 23.100 22.860 23.360 ;
        RECT 22.960 23.100 23.220 23.360 ;
        RECT 23.320 23.100 23.580 23.360 ;
        RECT 22.600 22.740 22.860 23.000 ;
        RECT 22.960 22.740 23.220 23.000 ;
        RECT 23.320 22.740 23.580 23.000 ;
        RECT 22.600 22.380 22.860 22.640 ;
        RECT 22.960 22.380 23.220 22.640 ;
        RECT 23.320 22.380 23.580 22.640 ;
        RECT 22.600 22.020 22.860 22.280 ;
        RECT 22.960 22.020 23.220 22.280 ;
        RECT 23.320 22.020 23.580 22.280 ;
        RECT 22.600 21.660 22.860 21.920 ;
        RECT 22.960 21.660 23.220 21.920 ;
        RECT 23.320 21.660 23.580 21.920 ;
        RECT 22.600 21.300 22.860 21.560 ;
        RECT 22.960 21.300 23.220 21.560 ;
        RECT 23.320 21.300 23.580 21.560 ;
        RECT 22.600 20.940 22.860 21.200 ;
        RECT 22.960 20.940 23.220 21.200 ;
        RECT 23.320 20.940 23.580 21.200 ;
        RECT 22.600 20.580 22.860 20.840 ;
        RECT 22.960 20.580 23.220 20.840 ;
        RECT 23.320 20.580 23.580 20.840 ;
        RECT 22.600 20.220 22.860 20.480 ;
        RECT 22.960 20.220 23.220 20.480 ;
        RECT 23.320 20.220 23.580 20.480 ;
        RECT 22.600 19.860 22.860 20.120 ;
        RECT 22.960 19.860 23.220 20.120 ;
        RECT 23.320 19.860 23.580 20.120 ;
        RECT 22.600 19.500 22.860 19.760 ;
        RECT 22.960 19.500 23.220 19.760 ;
        RECT 23.320 19.500 23.580 19.760 ;
        RECT 22.600 19.140 22.860 19.400 ;
        RECT 22.960 19.140 23.220 19.400 ;
        RECT 23.320 19.140 23.580 19.400 ;
        RECT 22.600 18.780 22.860 19.040 ;
        RECT 22.960 18.780 23.220 19.040 ;
        RECT 23.320 18.780 23.580 19.040 ;
        RECT 22.600 18.420 22.860 18.680 ;
        RECT 22.960 18.420 23.220 18.680 ;
        RECT 23.320 18.420 23.580 18.680 ;
        RECT 22.600 18.060 22.860 18.320 ;
        RECT 22.960 18.060 23.220 18.320 ;
        RECT 23.320 18.060 23.580 18.320 ;
        RECT 22.600 17.700 22.860 17.960 ;
        RECT 22.960 17.700 23.220 17.960 ;
        RECT 23.320 17.700 23.580 17.960 ;
        RECT 22.600 17.340 22.860 17.600 ;
        RECT 22.960 17.340 23.220 17.600 ;
        RECT 23.320 17.340 23.580 17.600 ;
        RECT 25.060 18.010 25.320 18.270 ;
        RECT 25.420 18.010 25.680 18.270 ;
        RECT 25.780 18.010 26.040 18.270 ;
        RECT 26.140 18.010 26.400 18.270 ;
        RECT 26.500 18.010 26.760 18.270 ;
        RECT 26.860 18.010 27.120 18.270 ;
        RECT 27.220 18.010 27.480 18.270 ;
        RECT 27.580 18.010 27.840 18.270 ;
        RECT 27.940 18.010 28.200 18.270 ;
        RECT 28.300 18.010 28.560 18.270 ;
        RECT 28.660 18.010 28.920 18.270 ;
        RECT 29.020 18.010 29.280 18.270 ;
        RECT 29.380 18.010 29.640 18.270 ;
        RECT 29.740 18.010 30.000 18.270 ;
        RECT 30.100 18.010 30.360 18.270 ;
        RECT 30.460 18.010 30.720 18.270 ;
        RECT 30.820 18.010 31.080 18.270 ;
        RECT 31.180 18.010 31.440 18.270 ;
        RECT 31.540 18.010 31.800 18.270 ;
        RECT 31.900 18.010 32.160 18.270 ;
        RECT 32.260 18.010 32.520 18.270 ;
        RECT 32.620 18.010 32.880 18.270 ;
        RECT 32.980 18.010 33.240 18.270 ;
        RECT 33.340 18.010 33.600 18.270 ;
        RECT 33.700 18.010 33.960 18.270 ;
        RECT 34.060 18.010 34.320 18.270 ;
        RECT 34.420 18.010 34.680 18.270 ;
        RECT 34.780 18.010 35.040 18.270 ;
        RECT 35.140 18.010 35.400 18.270 ;
        RECT 35.500 18.010 35.760 18.270 ;
        RECT 35.860 18.010 36.120 18.270 ;
        RECT 36.220 18.010 36.480 18.270 ;
        RECT 36.580 18.010 36.840 18.270 ;
        RECT 36.940 18.010 37.200 18.270 ;
        RECT 37.300 18.010 37.560 18.270 ;
        RECT 37.660 18.010 37.920 18.270 ;
        RECT 38.020 18.010 38.280 18.270 ;
        RECT 38.380 18.010 38.640 18.270 ;
        RECT 38.740 18.010 39.000 18.270 ;
        RECT 39.100 18.010 39.360 18.270 ;
        RECT 39.460 18.010 39.720 18.270 ;
        RECT 39.820 18.010 40.080 18.270 ;
        RECT 40.180 18.010 40.440 18.270 ;
        RECT 40.540 18.010 40.800 18.270 ;
        RECT 40.900 18.010 41.160 18.270 ;
        RECT 41.260 18.010 41.520 18.270 ;
        RECT 41.620 18.010 41.880 18.270 ;
        RECT 41.980 18.010 42.240 18.270 ;
        RECT 42.340 18.010 42.600 18.270 ;
        RECT 42.700 18.010 42.960 18.270 ;
        RECT 43.060 18.010 43.320 18.270 ;
        RECT 43.420 18.010 43.680 18.270 ;
        RECT 43.780 18.010 44.040 18.270 ;
        RECT 44.140 18.010 44.400 18.270 ;
        RECT 44.500 18.010 44.760 18.270 ;
        RECT 44.860 18.010 45.120 18.270 ;
        RECT 45.220 18.010 45.480 18.270 ;
        RECT 45.580 18.010 45.840 18.270 ;
        RECT 45.940 18.010 46.200 18.270 ;
        RECT 46.300 18.010 46.560 18.270 ;
        RECT 46.660 18.010 46.920 18.270 ;
        RECT 47.020 18.010 47.280 18.270 ;
        RECT 47.380 18.010 47.640 18.270 ;
        RECT 47.740 18.010 48.000 18.270 ;
        RECT 48.100 18.010 48.360 18.270 ;
        RECT 48.460 18.010 48.720 18.270 ;
        RECT 48.820 18.010 49.080 18.270 ;
        RECT 49.180 18.010 49.440 18.270 ;
        RECT 49.540 18.010 49.800 18.270 ;
        RECT 49.900 18.010 50.160 18.270 ;
        RECT 50.260 18.010 50.520 18.270 ;
        RECT 50.620 18.010 50.880 18.270 ;
        RECT 50.980 18.010 51.240 18.270 ;
        RECT 51.340 18.010 51.600 18.270 ;
        RECT 51.700 18.010 51.960 18.270 ;
        RECT 52.060 18.010 52.320 18.270 ;
        RECT 52.420 18.010 52.680 18.270 ;
        RECT 52.780 18.010 53.040 18.270 ;
        RECT 53.140 18.010 53.400 18.270 ;
        RECT 53.500 18.010 53.760 18.270 ;
        RECT 53.860 18.010 54.120 18.270 ;
        RECT 54.220 18.010 54.480 18.270 ;
        RECT 54.580 18.010 54.840 18.270 ;
        RECT 54.940 18.010 55.200 18.270 ;
        RECT 55.300 18.010 55.560 18.270 ;
        RECT 55.660 18.010 55.920 18.270 ;
        RECT 56.020 18.010 56.280 18.270 ;
        RECT 56.380 18.010 56.640 18.270 ;
        RECT 56.740 18.010 57.000 18.270 ;
        RECT 57.100 18.010 57.360 18.270 ;
        RECT 57.460 18.010 57.720 18.270 ;
        RECT 57.820 18.010 58.080 18.270 ;
        RECT 58.180 18.010 58.440 18.270 ;
        RECT 58.540 18.010 58.800 18.270 ;
        RECT 58.900 18.010 59.160 18.270 ;
        RECT 59.260 18.010 59.520 18.270 ;
        RECT 59.620 18.010 59.880 18.270 ;
        RECT 59.980 18.010 60.240 18.270 ;
        RECT 60.340 18.010 60.600 18.270 ;
        RECT 60.700 18.010 60.960 18.270 ;
        RECT 61.060 18.010 61.320 18.270 ;
        RECT 61.420 18.010 61.680 18.270 ;
        RECT 61.780 18.010 62.040 18.270 ;
        RECT 62.140 18.010 62.400 18.270 ;
        RECT 62.500 18.010 62.760 18.270 ;
        RECT 62.860 18.010 63.120 18.270 ;
        RECT 63.220 18.010 63.480 18.270 ;
        RECT 63.580 18.010 63.840 18.270 ;
        RECT 63.940 18.010 64.200 18.270 ;
        RECT 64.300 18.010 64.560 18.270 ;
        RECT 64.660 18.010 64.920 18.270 ;
        RECT 25.060 17.650 25.320 17.910 ;
        RECT 25.420 17.650 25.680 17.910 ;
        RECT 25.780 17.650 26.040 17.910 ;
        RECT 26.140 17.650 26.400 17.910 ;
        RECT 26.500 17.650 26.760 17.910 ;
        RECT 26.860 17.650 27.120 17.910 ;
        RECT 27.220 17.650 27.480 17.910 ;
        RECT 27.580 17.650 27.840 17.910 ;
        RECT 27.940 17.650 28.200 17.910 ;
        RECT 28.300 17.650 28.560 17.910 ;
        RECT 28.660 17.650 28.920 17.910 ;
        RECT 29.020 17.650 29.280 17.910 ;
        RECT 29.380 17.650 29.640 17.910 ;
        RECT 29.740 17.650 30.000 17.910 ;
        RECT 30.100 17.650 30.360 17.910 ;
        RECT 30.460 17.650 30.720 17.910 ;
        RECT 30.820 17.650 31.080 17.910 ;
        RECT 31.180 17.650 31.440 17.910 ;
        RECT 31.540 17.650 31.800 17.910 ;
        RECT 31.900 17.650 32.160 17.910 ;
        RECT 32.260 17.650 32.520 17.910 ;
        RECT 32.620 17.650 32.880 17.910 ;
        RECT 32.980 17.650 33.240 17.910 ;
        RECT 33.340 17.650 33.600 17.910 ;
        RECT 33.700 17.650 33.960 17.910 ;
        RECT 34.060 17.650 34.320 17.910 ;
        RECT 34.420 17.650 34.680 17.910 ;
        RECT 34.780 17.650 35.040 17.910 ;
        RECT 35.140 17.650 35.400 17.910 ;
        RECT 35.500 17.650 35.760 17.910 ;
        RECT 35.860 17.650 36.120 17.910 ;
        RECT 36.220 17.650 36.480 17.910 ;
        RECT 36.580 17.650 36.840 17.910 ;
        RECT 36.940 17.650 37.200 17.910 ;
        RECT 37.300 17.650 37.560 17.910 ;
        RECT 37.660 17.650 37.920 17.910 ;
        RECT 38.020 17.650 38.280 17.910 ;
        RECT 38.380 17.650 38.640 17.910 ;
        RECT 38.740 17.650 39.000 17.910 ;
        RECT 39.100 17.650 39.360 17.910 ;
        RECT 39.460 17.650 39.720 17.910 ;
        RECT 39.820 17.650 40.080 17.910 ;
        RECT 40.180 17.650 40.440 17.910 ;
        RECT 40.540 17.650 40.800 17.910 ;
        RECT 40.900 17.650 41.160 17.910 ;
        RECT 41.260 17.650 41.520 17.910 ;
        RECT 41.620 17.650 41.880 17.910 ;
        RECT 41.980 17.650 42.240 17.910 ;
        RECT 42.340 17.650 42.600 17.910 ;
        RECT 42.700 17.650 42.960 17.910 ;
        RECT 43.060 17.650 43.320 17.910 ;
        RECT 43.420 17.650 43.680 17.910 ;
        RECT 43.780 17.650 44.040 17.910 ;
        RECT 44.140 17.650 44.400 17.910 ;
        RECT 44.500 17.650 44.760 17.910 ;
        RECT 44.860 17.650 45.120 17.910 ;
        RECT 45.220 17.650 45.480 17.910 ;
        RECT 45.580 17.650 45.840 17.910 ;
        RECT 45.940 17.650 46.200 17.910 ;
        RECT 46.300 17.650 46.560 17.910 ;
        RECT 46.660 17.650 46.920 17.910 ;
        RECT 47.020 17.650 47.280 17.910 ;
        RECT 47.380 17.650 47.640 17.910 ;
        RECT 47.740 17.650 48.000 17.910 ;
        RECT 48.100 17.650 48.360 17.910 ;
        RECT 48.460 17.650 48.720 17.910 ;
        RECT 48.820 17.650 49.080 17.910 ;
        RECT 49.180 17.650 49.440 17.910 ;
        RECT 49.540 17.650 49.800 17.910 ;
        RECT 49.900 17.650 50.160 17.910 ;
        RECT 50.260 17.650 50.520 17.910 ;
        RECT 50.620 17.650 50.880 17.910 ;
        RECT 50.980 17.650 51.240 17.910 ;
        RECT 51.340 17.650 51.600 17.910 ;
        RECT 51.700 17.650 51.960 17.910 ;
        RECT 52.060 17.650 52.320 17.910 ;
        RECT 52.420 17.650 52.680 17.910 ;
        RECT 52.780 17.650 53.040 17.910 ;
        RECT 53.140 17.650 53.400 17.910 ;
        RECT 53.500 17.650 53.760 17.910 ;
        RECT 53.860 17.650 54.120 17.910 ;
        RECT 54.220 17.650 54.480 17.910 ;
        RECT 54.580 17.650 54.840 17.910 ;
        RECT 54.940 17.650 55.200 17.910 ;
        RECT 55.300 17.650 55.560 17.910 ;
        RECT 55.660 17.650 55.920 17.910 ;
        RECT 56.020 17.650 56.280 17.910 ;
        RECT 56.380 17.650 56.640 17.910 ;
        RECT 56.740 17.650 57.000 17.910 ;
        RECT 57.100 17.650 57.360 17.910 ;
        RECT 57.460 17.650 57.720 17.910 ;
        RECT 57.820 17.650 58.080 17.910 ;
        RECT 58.180 17.650 58.440 17.910 ;
        RECT 58.540 17.650 58.800 17.910 ;
        RECT 58.900 17.650 59.160 17.910 ;
        RECT 59.260 17.650 59.520 17.910 ;
        RECT 59.620 17.650 59.880 17.910 ;
        RECT 59.980 17.650 60.240 17.910 ;
        RECT 60.340 17.650 60.600 17.910 ;
        RECT 60.700 17.650 60.960 17.910 ;
        RECT 61.060 17.650 61.320 17.910 ;
        RECT 61.420 17.650 61.680 17.910 ;
        RECT 61.780 17.650 62.040 17.910 ;
        RECT 62.140 17.650 62.400 17.910 ;
        RECT 62.500 17.650 62.760 17.910 ;
        RECT 62.860 17.650 63.120 17.910 ;
        RECT 63.220 17.650 63.480 17.910 ;
        RECT 63.580 17.650 63.840 17.910 ;
        RECT 63.940 17.650 64.200 17.910 ;
        RECT 64.300 17.650 64.560 17.910 ;
        RECT 64.660 17.650 64.920 17.910 ;
        RECT 22.600 16.980 22.860 17.240 ;
        RECT 22.960 16.980 23.220 17.240 ;
        RECT 23.320 16.980 23.580 17.240 ;
        RECT 22.600 16.620 22.860 16.880 ;
        RECT 22.960 16.620 23.220 16.880 ;
        RECT 23.320 16.620 23.580 16.880 ;
        RECT 22.600 16.260 22.860 16.520 ;
        RECT 22.960 16.260 23.220 16.520 ;
        RECT 23.320 16.260 23.580 16.520 ;
        RECT 22.600 15.900 22.860 16.160 ;
        RECT 22.960 15.900 23.220 16.160 ;
        RECT 23.320 15.900 23.580 16.160 ;
        RECT 25.060 17.290 25.320 17.550 ;
        RECT 25.420 17.290 25.680 17.550 ;
        RECT 25.780 17.290 26.040 17.550 ;
        RECT 26.140 17.290 26.400 17.550 ;
        RECT 26.500 17.290 26.760 17.550 ;
        RECT 26.860 17.290 27.120 17.550 ;
        RECT 27.220 17.290 27.480 17.550 ;
        RECT 27.580 17.290 27.840 17.550 ;
        RECT 27.940 17.290 28.200 17.550 ;
        RECT 28.300 17.290 28.560 17.550 ;
        RECT 28.660 17.290 28.920 17.550 ;
        RECT 29.020 17.290 29.280 17.550 ;
        RECT 29.380 17.290 29.640 17.550 ;
        RECT 29.740 17.290 30.000 17.550 ;
        RECT 30.100 17.290 30.360 17.550 ;
        RECT 30.460 17.290 30.720 17.550 ;
        RECT 30.820 17.290 31.080 17.550 ;
        RECT 31.180 17.290 31.440 17.550 ;
        RECT 31.540 17.290 31.800 17.550 ;
        RECT 31.900 17.290 32.160 17.550 ;
        RECT 32.260 17.290 32.520 17.550 ;
        RECT 32.620 17.290 32.880 17.550 ;
        RECT 32.980 17.290 33.240 17.550 ;
        RECT 33.340 17.290 33.600 17.550 ;
        RECT 33.700 17.290 33.960 17.550 ;
        RECT 34.060 17.290 34.320 17.550 ;
        RECT 34.420 17.290 34.680 17.550 ;
        RECT 34.780 17.290 35.040 17.550 ;
        RECT 35.140 17.290 35.400 17.550 ;
        RECT 35.500 17.290 35.760 17.550 ;
        RECT 35.860 17.290 36.120 17.550 ;
        RECT 36.220 17.290 36.480 17.550 ;
        RECT 36.580 17.290 36.840 17.550 ;
        RECT 36.940 17.290 37.200 17.550 ;
        RECT 37.300 17.290 37.560 17.550 ;
        RECT 37.660 17.290 37.920 17.550 ;
        RECT 38.020 17.290 38.280 17.550 ;
        RECT 38.380 17.290 38.640 17.550 ;
        RECT 38.740 17.290 39.000 17.550 ;
        RECT 39.100 17.290 39.360 17.550 ;
        RECT 39.460 17.290 39.720 17.550 ;
        RECT 39.820 17.290 40.080 17.550 ;
        RECT 40.180 17.290 40.440 17.550 ;
        RECT 40.540 17.290 40.800 17.550 ;
        RECT 40.900 17.290 41.160 17.550 ;
        RECT 41.260 17.290 41.520 17.550 ;
        RECT 41.620 17.290 41.880 17.550 ;
        RECT 41.980 17.290 42.240 17.550 ;
        RECT 42.340 17.290 42.600 17.550 ;
        RECT 42.700 17.290 42.960 17.550 ;
        RECT 43.060 17.290 43.320 17.550 ;
        RECT 43.420 17.290 43.680 17.550 ;
        RECT 43.780 17.290 44.040 17.550 ;
        RECT 44.140 17.290 44.400 17.550 ;
        RECT 44.500 17.290 44.760 17.550 ;
        RECT 44.860 17.290 45.120 17.550 ;
        RECT 45.220 17.290 45.480 17.550 ;
        RECT 45.580 17.290 45.840 17.550 ;
        RECT 45.940 17.290 46.200 17.550 ;
        RECT 46.300 17.290 46.560 17.550 ;
        RECT 46.660 17.290 46.920 17.550 ;
        RECT 47.020 17.290 47.280 17.550 ;
        RECT 47.380 17.290 47.640 17.550 ;
        RECT 47.740 17.290 48.000 17.550 ;
        RECT 48.100 17.290 48.360 17.550 ;
        RECT 48.460 17.290 48.720 17.550 ;
        RECT 48.820 17.290 49.080 17.550 ;
        RECT 49.180 17.290 49.440 17.550 ;
        RECT 49.540 17.290 49.800 17.550 ;
        RECT 49.900 17.290 50.160 17.550 ;
        RECT 50.260 17.290 50.520 17.550 ;
        RECT 50.620 17.290 50.880 17.550 ;
        RECT 50.980 17.290 51.240 17.550 ;
        RECT 51.340 17.290 51.600 17.550 ;
        RECT 51.700 17.290 51.960 17.550 ;
        RECT 52.060 17.290 52.320 17.550 ;
        RECT 52.420 17.290 52.680 17.550 ;
        RECT 52.780 17.290 53.040 17.550 ;
        RECT 53.140 17.290 53.400 17.550 ;
        RECT 53.500 17.290 53.760 17.550 ;
        RECT 53.860 17.290 54.120 17.550 ;
        RECT 54.220 17.290 54.480 17.550 ;
        RECT 54.580 17.290 54.840 17.550 ;
        RECT 54.940 17.290 55.200 17.550 ;
        RECT 55.300 17.290 55.560 17.550 ;
        RECT 55.660 17.290 55.920 17.550 ;
        RECT 56.020 17.290 56.280 17.550 ;
        RECT 56.380 17.290 56.640 17.550 ;
        RECT 56.740 17.290 57.000 17.550 ;
        RECT 57.100 17.290 57.360 17.550 ;
        RECT 57.460 17.290 57.720 17.550 ;
        RECT 57.820 17.290 58.080 17.550 ;
        RECT 58.180 17.290 58.440 17.550 ;
        RECT 58.540 17.290 58.800 17.550 ;
        RECT 58.900 17.290 59.160 17.550 ;
        RECT 59.260 17.290 59.520 17.550 ;
        RECT 59.620 17.290 59.880 17.550 ;
        RECT 59.980 17.290 60.240 17.550 ;
        RECT 60.340 17.290 60.600 17.550 ;
        RECT 60.700 17.290 60.960 17.550 ;
        RECT 61.060 17.290 61.320 17.550 ;
        RECT 61.420 17.290 61.680 17.550 ;
        RECT 61.780 17.290 62.040 17.550 ;
        RECT 62.140 17.290 62.400 17.550 ;
        RECT 62.500 17.290 62.760 17.550 ;
        RECT 62.860 17.290 63.120 17.550 ;
        RECT 63.220 17.290 63.480 17.550 ;
        RECT 63.580 17.290 63.840 17.550 ;
        RECT 63.940 17.290 64.200 17.550 ;
        RECT 64.300 17.290 64.560 17.550 ;
        RECT 64.660 17.290 64.920 17.550 ;
        RECT 22.600 15.540 22.860 15.800 ;
        RECT 22.960 15.540 23.220 15.800 ;
        RECT 23.320 15.540 23.580 15.800 ;
        RECT 22.600 15.180 22.860 15.440 ;
        RECT 22.960 15.180 23.220 15.440 ;
        RECT 23.320 15.180 23.580 15.440 ;
        RECT 22.600 14.820 22.860 15.080 ;
        RECT 22.960 14.820 23.220 15.080 ;
        RECT 23.320 14.820 23.580 15.080 ;
        RECT 22.600 14.460 22.860 14.720 ;
        RECT 22.960 14.460 23.220 14.720 ;
        RECT 23.320 14.460 23.580 14.720 ;
        RECT 22.600 14.100 22.860 14.360 ;
        RECT 22.960 14.100 23.220 14.360 ;
        RECT 23.320 14.100 23.580 14.360 ;
        RECT 22.600 13.740 22.860 14.000 ;
        RECT 22.960 13.740 23.220 14.000 ;
        RECT 23.320 13.740 23.580 14.000 ;
        RECT 22.600 13.380 22.860 13.640 ;
        RECT 22.960 13.380 23.220 13.640 ;
        RECT 23.320 13.380 23.580 13.640 ;
        RECT 22.600 13.020 22.860 13.280 ;
        RECT 22.960 13.020 23.220 13.280 ;
        RECT 23.320 13.020 23.580 13.280 ;
        RECT 22.600 12.660 22.860 12.920 ;
        RECT 22.960 12.660 23.220 12.920 ;
        RECT 23.320 12.660 23.580 12.920 ;
        RECT 22.600 12.300 22.860 12.560 ;
        RECT 22.960 12.300 23.220 12.560 ;
        RECT 23.320 12.300 23.580 12.560 ;
        RECT 22.600 11.940 22.860 12.200 ;
        RECT 22.960 11.940 23.220 12.200 ;
        RECT 23.320 11.940 23.580 12.200 ;
        RECT 22.600 11.580 22.860 11.840 ;
        RECT 22.960 11.580 23.220 11.840 ;
        RECT 23.320 11.580 23.580 11.840 ;
        RECT 22.600 11.220 22.860 11.480 ;
        RECT 22.960 11.220 23.220 11.480 ;
        RECT 23.320 11.220 23.580 11.480 ;
        RECT 22.600 10.860 22.860 11.120 ;
        RECT 22.960 10.860 23.220 11.120 ;
        RECT 23.320 10.860 23.580 11.120 ;
        RECT 22.600 10.500 22.860 10.760 ;
        RECT 22.960 10.500 23.220 10.760 ;
        RECT 23.320 10.500 23.580 10.760 ;
        RECT 22.600 10.140 22.860 10.400 ;
        RECT 22.960 10.140 23.220 10.400 ;
        RECT 23.320 10.140 23.580 10.400 ;
        RECT 22.600 9.780 22.860 10.040 ;
        RECT 22.960 9.780 23.220 10.040 ;
        RECT 23.320 9.780 23.580 10.040 ;
        RECT 22.600 9.420 22.860 9.680 ;
        RECT 22.960 9.420 23.220 9.680 ;
        RECT 23.320 9.420 23.580 9.680 ;
        RECT 22.600 9.060 22.860 9.320 ;
        RECT 22.960 9.060 23.220 9.320 ;
        RECT 23.320 9.060 23.580 9.320 ;
        RECT 22.600 8.700 22.860 8.960 ;
        RECT 22.960 8.700 23.220 8.960 ;
        RECT 23.320 8.700 23.580 8.960 ;
        RECT 22.600 8.340 22.860 8.600 ;
        RECT 22.960 8.340 23.220 8.600 ;
        RECT 23.320 8.340 23.580 8.600 ;
        RECT 22.600 7.980 22.860 8.240 ;
        RECT 22.960 7.980 23.220 8.240 ;
        RECT 23.320 7.980 23.580 8.240 ;
        RECT 22.600 7.620 22.860 7.880 ;
        RECT 22.960 7.620 23.220 7.880 ;
        RECT 23.320 7.620 23.580 7.880 ;
        RECT 22.600 7.260 22.860 7.520 ;
        RECT 22.960 7.260 23.220 7.520 ;
        RECT 23.320 7.260 23.580 7.520 ;
        RECT 22.600 6.900 22.860 7.160 ;
        RECT 22.960 6.900 23.220 7.160 ;
        RECT 23.320 6.900 23.580 7.160 ;
      LAYER met2 ;
        RECT 21.430 108.930 21.810 110.425 ;
        RECT 24.190 108.930 24.570 110.425 ;
        RECT 26.950 108.930 27.330 110.425 ;
        RECT 29.710 108.930 30.090 110.425 ;
        RECT 32.470 108.930 32.850 110.425 ;
        RECT 35.230 108.930 35.610 110.425 ;
        RECT 37.990 108.930 38.370 110.425 ;
        RECT 40.750 108.930 41.130 110.425 ;
        RECT 85.455 103.480 102.475 103.960 ;
        RECT 107.185 101.980 109.355 102.350 ;
        RECT 11.610 90.805 51.530 91.845 ;
        RECT 56.820 88.905 96.740 89.945 ;
        RECT 16.520 47.970 17.560 87.890 ;
        RECT 99.195 49.300 100.235 89.220 ;
        RECT 22.570 6.870 23.610 46.790 ;
        RECT 65.225 26.855 105.145 27.895 ;
        RECT 25.030 17.260 64.950 18.300 ;
      LAYER via2 ;
        RECT 21.480 110.100 21.760 110.380 ;
        RECT 21.480 109.700 21.760 109.980 ;
        RECT 24.240 110.100 24.520 110.380 ;
        RECT 24.240 109.700 24.520 109.980 ;
        RECT 27.000 110.100 27.280 110.380 ;
        RECT 27.000 109.700 27.280 109.980 ;
        RECT 29.760 110.100 30.040 110.380 ;
        RECT 29.760 109.700 30.040 109.980 ;
        RECT 32.520 110.100 32.800 110.380 ;
        RECT 32.520 109.700 32.800 109.980 ;
        RECT 35.280 110.100 35.560 110.380 ;
        RECT 35.280 109.700 35.560 109.980 ;
        RECT 38.040 110.100 38.320 110.380 ;
        RECT 38.040 109.700 38.320 109.980 ;
        RECT 40.800 110.100 41.080 110.380 ;
        RECT 40.800 109.700 41.080 109.980 ;
        RECT 85.625 103.580 85.905 103.860 ;
        RECT 86.025 103.580 86.305 103.860 ;
        RECT 86.425 103.580 86.705 103.860 ;
        RECT 86.825 103.580 87.105 103.860 ;
        RECT 87.225 103.580 87.505 103.860 ;
        RECT 87.625 103.580 87.905 103.860 ;
        RECT 88.025 103.580 88.305 103.860 ;
        RECT 88.425 103.580 88.705 103.860 ;
        RECT 88.825 103.580 89.105 103.860 ;
        RECT 89.225 103.580 89.505 103.860 ;
        RECT 89.625 103.580 89.905 103.860 ;
        RECT 90.025 103.580 90.305 103.860 ;
        RECT 90.425 103.580 90.705 103.860 ;
        RECT 90.825 103.580 91.105 103.860 ;
        RECT 91.225 103.580 91.505 103.860 ;
        RECT 91.625 103.580 91.905 103.860 ;
        RECT 92.025 103.580 92.305 103.860 ;
        RECT 92.425 103.580 92.705 103.860 ;
        RECT 92.825 103.580 93.105 103.860 ;
        RECT 93.225 103.580 93.505 103.860 ;
        RECT 93.625 103.580 93.905 103.860 ;
        RECT 94.025 103.580 94.305 103.860 ;
        RECT 94.425 103.580 94.705 103.860 ;
        RECT 94.825 103.580 95.105 103.860 ;
        RECT 95.225 103.580 95.505 103.860 ;
        RECT 95.625 103.580 95.905 103.860 ;
        RECT 96.025 103.580 96.305 103.860 ;
        RECT 96.425 103.580 96.705 103.860 ;
        RECT 96.825 103.580 97.105 103.860 ;
        RECT 97.225 103.580 97.505 103.860 ;
        RECT 97.625 103.580 97.905 103.860 ;
        RECT 98.025 103.580 98.305 103.860 ;
        RECT 98.425 103.580 98.705 103.860 ;
        RECT 98.825 103.580 99.105 103.860 ;
        RECT 99.225 103.580 99.505 103.860 ;
        RECT 99.625 103.580 99.905 103.860 ;
        RECT 100.025 103.580 100.305 103.860 ;
        RECT 100.425 103.580 100.705 103.860 ;
        RECT 100.825 103.580 101.105 103.860 ;
        RECT 101.225 103.580 101.505 103.860 ;
        RECT 101.625 103.580 101.905 103.860 ;
        RECT 102.025 103.580 102.305 103.860 ;
        RECT 107.230 102.025 107.510 102.305 ;
        RECT 107.680 102.025 107.960 102.305 ;
        RECT 108.130 102.025 108.410 102.305 ;
        RECT 108.580 102.025 108.860 102.305 ;
        RECT 109.030 102.025 109.310 102.305 ;
        RECT 11.830 90.985 51.310 91.665 ;
        RECT 57.040 89.085 96.520 89.765 ;
        RECT 16.700 48.190 17.380 87.670 ;
        RECT 99.375 49.520 100.055 89.000 ;
        RECT 22.750 7.090 23.430 46.570 ;
        RECT 65.445 27.030 104.925 27.710 ;
        RECT 25.250 17.440 64.730 18.120 ;
      LAYER met3 ;
        RECT 0.000 106.850 41.130 111.520 ;
        RECT 139.580 106.850 153.165 111.520 ;
        RECT 0.000 0.000 153.165 106.850 ;
      LAYER via3 ;
        RECT 0.240 0.200 1.760 111.320 ;
        RECT 21.460 110.880 21.780 111.200 ;
        RECT 24.220 110.880 24.540 111.200 ;
        RECT 26.980 110.880 27.300 111.200 ;
        RECT 29.740 110.880 30.060 111.200 ;
        RECT 32.500 110.880 32.820 111.200 ;
        RECT 35.260 110.880 35.580 111.200 ;
        RECT 38.020 110.880 38.340 111.200 ;
        RECT 40.780 110.880 41.100 111.200 ;
        RECT 21.460 110.480 21.780 110.800 ;
        RECT 24.220 110.480 24.540 110.800 ;
        RECT 26.980 110.480 27.300 110.800 ;
        RECT 29.740 110.480 30.060 110.800 ;
        RECT 32.500 110.480 32.820 110.800 ;
        RECT 35.260 110.480 35.580 110.800 ;
        RECT 38.020 110.480 38.340 110.800 ;
        RECT 40.780 110.480 41.100 110.800 ;
      LAYER met4 ;
        RECT 0.000 0.000 2.000 111.520 ;
        RECT 21.470 111.230 21.770 111.520 ;
        RECT 24.230 111.230 24.530 111.520 ;
        RECT 26.990 111.230 27.290 111.520 ;
        RECT 29.750 111.230 30.050 111.520 ;
        RECT 32.510 111.230 32.810 111.520 ;
        RECT 35.270 111.230 35.570 111.520 ;
        RECT 38.030 111.230 38.330 111.520 ;
        RECT 40.790 111.230 41.090 111.520 ;
        RECT 21.430 110.450 21.810 111.230 ;
        RECT 24.190 110.450 24.570 111.230 ;
        RECT 26.950 110.450 27.330 111.230 ;
        RECT 29.710 110.450 30.090 111.230 ;
        RECT 32.470 110.450 32.850 111.230 ;
        RECT 35.230 110.450 35.610 111.230 ;
        RECT 37.990 110.450 38.370 111.230 ;
        RECT 40.750 110.450 41.130 111.230 ;
    END
  END uio_oe[0]
  PIN uo_out[0]
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER li1 ;
        RECT 90.610 106.180 90.780 106.185 ;
        RECT 91.450 106.180 91.620 106.185 ;
        RECT 92.290 106.180 92.540 106.185 ;
        RECT 85.540 105.705 85.815 106.075 ;
        RECT 86.330 105.705 86.660 106.180 ;
        RECT 87.170 105.705 87.500 106.180 ;
        RECT 88.010 105.705 88.340 106.180 ;
        RECT 88.850 105.705 89.180 106.180 ;
        RECT 89.690 105.705 90.020 106.180 ;
        RECT 90.530 105.705 90.860 106.180 ;
        RECT 91.370 105.705 91.700 106.180 ;
        RECT 92.210 105.705 92.540 106.180 ;
        RECT 85.540 105.535 92.540 105.705 ;
        RECT 85.540 104.995 85.920 105.535 ;
        RECT 85.540 104.825 92.540 104.995 ;
        RECT 85.540 104.080 85.815 104.825 ;
        RECT 86.330 103.975 86.660 104.825 ;
        RECT 87.170 103.975 87.500 104.825 ;
        RECT 88.010 103.975 88.340 104.825 ;
        RECT 88.850 103.975 89.180 104.825 ;
        RECT 89.690 103.975 90.020 104.825 ;
        RECT 90.530 103.975 90.860 104.825 ;
        RECT 91.370 103.975 91.700 104.825 ;
        RECT 92.210 103.975 92.540 104.825 ;
      LAYER mcon ;
        RECT 85.590 105.860 85.760 106.030 ;
        RECT 85.590 105.430 85.760 105.600 ;
        RECT 85.590 104.995 85.760 105.165 ;
        RECT 85.590 104.560 85.760 104.730 ;
        RECT 85.590 104.130 85.760 104.300 ;
      LAYER met1 ;
        RECT 84.915 106.060 85.285 109.650 ;
        RECT 84.915 104.100 85.815 106.060 ;
      LAYER via ;
        RECT 84.970 109.335 85.230 109.595 ;
        RECT 84.970 108.985 85.230 109.245 ;
      LAYER met2 ;
        RECT 84.910 108.930 85.290 110.425 ;
      LAYER via2 ;
        RECT 84.960 110.100 85.240 110.380 ;
        RECT 84.960 109.700 85.240 109.980 ;
      LAYER met3 ;
        RECT 84.910 109.650 85.290 111.230 ;
      LAYER via3 ;
        RECT 84.940 110.880 85.260 111.200 ;
        RECT 84.940 110.480 85.260 110.800 ;
      LAYER met4 ;
        RECT 84.950 111.230 85.250 111.520 ;
        RECT 84.910 110.450 85.290 111.230 ;
    END
  END uo_out[0]
  OBS
      LAYER pwell ;
        RECT 95.255 106.335 95.425 106.525 ;
        RECT 100.775 106.335 100.945 106.525 ;
        RECT 102.150 106.335 102.320 106.525 ;
        RECT 85.820 105.425 95.570 106.335 ;
        RECT 95.960 105.425 101.090 106.335 ;
        RECT 101.100 105.555 102.470 106.335 ;
      LAYER nwell ;
        RECT 85.265 103.530 102.665 105.135 ;
      LAYER li1 ;
        RECT 117.035 107.070 119.215 107.420 ;
        RECT 119.615 107.070 121.795 107.420 ;
        RECT 93.050 105.705 93.380 106.180 ;
        RECT 93.890 105.705 94.220 106.180 ;
        RECT 94.730 105.705 95.060 106.180 ;
        RECT 92.710 105.535 95.060 105.705 ;
        RECT 96.550 105.705 96.720 106.185 ;
        RECT 97.390 105.705 97.560 106.185 ;
        RECT 98.230 105.705 98.400 106.185 ;
        RECT 99.070 105.705 99.240 106.185 ;
        RECT 99.910 105.705 100.080 106.180 ;
        RECT 100.750 105.705 100.920 106.185 ;
        RECT 96.550 105.535 99.240 105.705 ;
        RECT 99.500 105.535 100.920 105.705 ;
        RECT 101.180 105.680 101.440 106.185 ;
        RECT 102.130 105.805 102.300 106.185 ;
        RECT 92.710 105.365 92.885 105.535 ;
        RECT 96.550 105.365 96.805 105.535 ;
        RECT 99.500 105.365 99.675 105.535 ;
        RECT 101.180 105.365 101.360 105.680 ;
        RECT 101.635 105.635 102.300 105.805 ;
        RECT 114.550 105.800 116.730 106.150 ;
        RECT 122.100 105.800 124.280 106.150 ;
        RECT 101.635 105.380 101.805 105.635 ;
        RECT 86.165 105.165 92.885 105.365 ;
        RECT 93.090 105.165 96.805 105.365 ;
        RECT 97.050 105.195 99.675 105.365 ;
        RECT 92.710 104.995 92.885 105.165 ;
        RECT 96.550 104.995 96.805 105.165 ;
        RECT 99.500 104.995 99.675 105.195 ;
        RECT 99.855 105.165 101.360 105.365 ;
        RECT 92.710 104.825 95.060 104.995 ;
        RECT 93.050 103.975 93.380 104.825 ;
        RECT 93.890 103.975 94.220 104.825 ;
        RECT 94.730 103.975 95.060 104.825 ;
        RECT 96.550 104.825 99.240 104.995 ;
        RECT 99.500 104.825 101.000 104.995 ;
        RECT 96.550 103.975 96.720 104.825 ;
        RECT 97.390 103.975 97.560 104.825 ;
        RECT 98.230 103.975 98.400 104.825 ;
        RECT 99.070 103.975 99.240 104.825 ;
        RECT 99.830 103.975 100.160 104.825 ;
        RECT 100.670 103.975 101.000 104.825 ;
        RECT 101.180 104.880 101.360 105.165 ;
        RECT 101.530 105.050 101.805 105.380 ;
        RECT 102.030 105.085 102.690 105.455 ;
        RECT 101.635 104.905 101.805 105.050 ;
        RECT 101.180 103.975 101.450 104.880 ;
        RECT 101.635 104.735 102.310 104.905 ;
        RECT 102.130 103.975 102.310 104.735 ;
        RECT 112.065 104.530 114.245 104.880 ;
        RECT 124.585 104.530 126.765 104.880 ;
        RECT 109.580 103.260 111.760 103.610 ;
        RECT 127.070 103.260 129.250 103.610 ;
        RECT 11.040 102.175 11.210 102.505 ;
        RECT 11.645 102.005 12.335 102.175 ;
        RECT 109.575 101.985 111.765 102.345 ;
        RECT 112.155 101.985 114.345 102.345 ;
        RECT 114.545 101.985 116.735 102.345 ;
        RECT 117.125 101.985 119.315 102.345 ;
        RECT 119.515 101.985 121.705 102.345 ;
        RECT 122.095 101.985 124.285 102.345 ;
        RECT 124.485 101.985 126.675 102.345 ;
        RECT 127.070 101.990 129.250 102.340 ;
        RECT 11.645 101.185 41.495 101.715 ;
        RECT 11.120 99.235 11.290 101.005 ;
        RECT 109.670 100.715 111.860 101.075 ;
        RECT 112.060 100.715 114.250 101.075 ;
        RECT 114.640 100.715 116.830 101.075 ;
        RECT 117.030 100.715 119.220 101.075 ;
        RECT 119.610 100.715 121.800 101.075 ;
        RECT 122.000 100.715 124.190 101.075 ;
        RECT 124.580 100.715 126.770 101.075 ;
        RECT 126.970 100.715 129.160 101.075 ;
        RECT 56.250 100.275 56.420 100.605 ;
        RECT 56.855 100.105 57.545 100.275 ;
        RECT 56.855 99.285 86.705 99.815 ;
        RECT 11.645 98.525 41.495 99.055 ;
        RECT 11.605 97.075 51.535 97.965 ;
        RECT 56.330 97.335 56.500 99.105 ;
        RECT 11.120 93.045 11.290 96.975 ;
        RECT 56.855 96.625 86.705 97.155 ;
        RECT 56.815 95.175 96.745 96.065 ;
        RECT 56.330 91.145 56.500 95.075 ;
        RECT 101.435 89.540 105.365 89.710 ;
        RECT 107.625 89.540 109.395 89.710 ;
        RECT 110.565 89.620 110.895 89.790 ;
        RECT 6.190 48.005 6.360 48.695 ;
        RECT 6.650 48.005 7.180 77.855 ;
        RECT 9.310 48.005 9.840 77.855 ;
        RECT 10.400 47.965 11.290 87.895 ;
        RECT 105.465 49.295 106.355 89.225 ;
        RECT 106.915 59.335 107.445 89.185 ;
        RECT 109.575 59.335 110.105 89.185 ;
        RECT 110.395 88.495 110.565 89.185 ;
        RECT 5.860 47.400 6.190 47.570 ;
        RECT 7.360 47.480 9.130 47.650 ;
        RECT 11.390 47.480 15.320 47.650 ;
        RECT 12.240 6.905 12.410 7.595 ;
        RECT 12.700 6.905 13.230 36.755 ;
        RECT 15.360 6.905 15.890 36.755 ;
        RECT 16.450 6.865 17.340 46.795 ;
        RECT 105.465 21.725 105.635 25.655 ;
        RECT 65.220 20.735 105.150 21.625 ;
        RECT 75.260 19.645 105.110 20.175 ;
        RECT 105.465 17.695 105.635 19.465 ;
        RECT 75.260 16.985 105.110 17.515 ;
        RECT 104.420 16.525 105.110 16.695 ;
        RECT 105.545 16.195 105.715 16.525 ;
        RECT 65.270 12.130 65.440 16.060 ;
        RECT 25.025 11.140 64.955 12.030 ;
        RECT 35.065 10.050 64.915 10.580 ;
        RECT 65.270 8.100 65.440 9.870 ;
        RECT 35.065 7.390 64.915 7.920 ;
        RECT 64.225 6.930 64.915 7.100 ;
        RECT 65.350 6.600 65.520 6.930 ;
        RECT 11.910 6.300 12.240 6.470 ;
        RECT 13.410 6.380 15.180 6.550 ;
        RECT 17.440 6.380 21.370 6.550 ;
      LAYER mcon ;
        RECT 117.145 107.160 117.315 107.330 ;
        RECT 117.505 107.160 117.675 107.330 ;
        RECT 117.865 107.160 118.035 107.330 ;
        RECT 118.225 107.160 118.395 107.330 ;
        RECT 118.585 107.160 118.755 107.330 ;
        RECT 118.945 107.160 119.115 107.330 ;
        RECT 119.710 107.160 119.880 107.330 ;
        RECT 120.070 107.160 120.240 107.330 ;
        RECT 120.430 107.160 120.600 107.330 ;
        RECT 120.790 107.160 120.960 107.330 ;
        RECT 121.150 107.160 121.320 107.330 ;
        RECT 121.510 107.160 121.680 107.330 ;
        RECT 114.660 105.890 114.830 106.060 ;
        RECT 115.020 105.890 115.190 106.060 ;
        RECT 115.380 105.890 115.550 106.060 ;
        RECT 115.740 105.890 115.910 106.060 ;
        RECT 116.100 105.890 116.270 106.060 ;
        RECT 116.460 105.890 116.630 106.060 ;
        RECT 122.195 105.890 122.365 106.060 ;
        RECT 122.555 105.890 122.725 106.060 ;
        RECT 122.915 105.890 123.085 106.060 ;
        RECT 123.275 105.890 123.445 106.060 ;
        RECT 123.635 105.890 123.805 106.060 ;
        RECT 123.995 105.890 124.165 106.060 ;
        RECT 102.085 105.180 102.255 105.350 ;
        RECT 102.480 105.180 102.650 105.350 ;
        RECT 112.175 104.620 112.345 104.790 ;
        RECT 112.535 104.620 112.705 104.790 ;
        RECT 112.895 104.620 113.065 104.790 ;
        RECT 113.255 104.620 113.425 104.790 ;
        RECT 113.615 104.620 113.785 104.790 ;
        RECT 113.975 104.620 114.145 104.790 ;
        RECT 124.680 104.620 124.850 104.790 ;
        RECT 125.040 104.620 125.210 104.790 ;
        RECT 125.400 104.620 125.570 104.790 ;
        RECT 125.760 104.620 125.930 104.790 ;
        RECT 126.120 104.620 126.290 104.790 ;
        RECT 126.480 104.620 126.650 104.790 ;
        RECT 109.690 103.350 109.860 103.520 ;
        RECT 110.050 103.350 110.220 103.520 ;
        RECT 110.410 103.350 110.580 103.520 ;
        RECT 110.770 103.350 110.940 103.520 ;
        RECT 111.130 103.350 111.300 103.520 ;
        RECT 111.490 103.350 111.660 103.520 ;
        RECT 127.165 103.350 127.335 103.520 ;
        RECT 127.525 103.350 127.695 103.520 ;
        RECT 127.885 103.350 128.055 103.520 ;
        RECT 128.245 103.350 128.415 103.520 ;
        RECT 128.605 103.350 128.775 103.520 ;
        RECT 128.965 103.350 129.135 103.520 ;
        RECT 11.040 102.255 11.210 102.425 ;
        RECT 11.725 102.005 11.895 102.175 ;
        RECT 12.085 102.005 12.255 102.175 ;
        RECT 109.690 102.080 109.860 102.250 ;
        RECT 110.050 102.080 110.220 102.250 ;
        RECT 110.410 102.080 110.580 102.250 ;
        RECT 110.770 102.080 110.940 102.250 ;
        RECT 111.130 102.080 111.300 102.250 ;
        RECT 111.490 102.080 111.660 102.250 ;
        RECT 112.255 102.080 112.425 102.250 ;
        RECT 112.615 102.080 112.785 102.250 ;
        RECT 112.975 102.080 113.145 102.250 ;
        RECT 113.335 102.080 113.505 102.250 ;
        RECT 113.695 102.080 113.865 102.250 ;
        RECT 114.055 102.080 114.225 102.250 ;
        RECT 114.660 102.080 114.830 102.250 ;
        RECT 115.020 102.080 115.190 102.250 ;
        RECT 115.380 102.080 115.550 102.250 ;
        RECT 115.740 102.080 115.910 102.250 ;
        RECT 116.100 102.080 116.270 102.250 ;
        RECT 116.460 102.080 116.630 102.250 ;
        RECT 117.225 102.080 117.395 102.250 ;
        RECT 117.585 102.080 117.755 102.250 ;
        RECT 117.945 102.080 118.115 102.250 ;
        RECT 118.305 102.080 118.475 102.250 ;
        RECT 118.665 102.080 118.835 102.250 ;
        RECT 119.025 102.080 119.195 102.250 ;
        RECT 119.630 102.080 119.800 102.250 ;
        RECT 119.990 102.080 120.160 102.250 ;
        RECT 120.350 102.080 120.520 102.250 ;
        RECT 120.710 102.080 120.880 102.250 ;
        RECT 121.070 102.080 121.240 102.250 ;
        RECT 121.430 102.080 121.600 102.250 ;
        RECT 122.195 102.080 122.365 102.250 ;
        RECT 122.555 102.080 122.725 102.250 ;
        RECT 122.915 102.080 123.085 102.250 ;
        RECT 123.275 102.080 123.445 102.250 ;
        RECT 123.635 102.080 123.805 102.250 ;
        RECT 123.995 102.080 124.165 102.250 ;
        RECT 124.600 102.080 124.770 102.250 ;
        RECT 124.960 102.080 125.130 102.250 ;
        RECT 125.320 102.080 125.490 102.250 ;
        RECT 125.680 102.080 125.850 102.250 ;
        RECT 126.040 102.080 126.210 102.250 ;
        RECT 126.400 102.080 126.570 102.250 ;
        RECT 127.165 102.080 127.335 102.250 ;
        RECT 127.525 102.080 127.695 102.250 ;
        RECT 127.885 102.080 128.055 102.250 ;
        RECT 128.245 102.080 128.415 102.250 ;
        RECT 128.605 102.080 128.775 102.250 ;
        RECT 128.965 102.080 129.135 102.250 ;
        RECT 11.725 101.185 41.415 101.715 ;
        RECT 11.120 100.755 11.290 100.925 ;
        RECT 109.770 100.810 109.940 100.980 ;
        RECT 110.130 100.810 110.300 100.980 ;
        RECT 110.490 100.810 110.660 100.980 ;
        RECT 110.850 100.810 111.020 100.980 ;
        RECT 111.210 100.810 111.380 100.980 ;
        RECT 111.570 100.810 111.740 100.980 ;
        RECT 112.175 100.810 112.345 100.980 ;
        RECT 112.535 100.810 112.705 100.980 ;
        RECT 112.895 100.810 113.065 100.980 ;
        RECT 113.255 100.810 113.425 100.980 ;
        RECT 113.615 100.810 113.785 100.980 ;
        RECT 113.975 100.810 114.145 100.980 ;
        RECT 114.740 100.810 114.910 100.980 ;
        RECT 115.100 100.810 115.270 100.980 ;
        RECT 115.460 100.810 115.630 100.980 ;
        RECT 115.820 100.810 115.990 100.980 ;
        RECT 116.180 100.810 116.350 100.980 ;
        RECT 116.540 100.810 116.710 100.980 ;
        RECT 117.145 100.810 117.315 100.980 ;
        RECT 117.505 100.810 117.675 100.980 ;
        RECT 117.865 100.810 118.035 100.980 ;
        RECT 118.225 100.810 118.395 100.980 ;
        RECT 118.585 100.810 118.755 100.980 ;
        RECT 118.945 100.810 119.115 100.980 ;
        RECT 119.710 100.810 119.880 100.980 ;
        RECT 120.070 100.810 120.240 100.980 ;
        RECT 120.430 100.810 120.600 100.980 ;
        RECT 120.790 100.810 120.960 100.980 ;
        RECT 121.150 100.810 121.320 100.980 ;
        RECT 121.510 100.810 121.680 100.980 ;
        RECT 122.115 100.810 122.285 100.980 ;
        RECT 122.475 100.810 122.645 100.980 ;
        RECT 122.835 100.810 123.005 100.980 ;
        RECT 123.195 100.810 123.365 100.980 ;
        RECT 123.555 100.810 123.725 100.980 ;
        RECT 123.915 100.810 124.085 100.980 ;
        RECT 124.680 100.810 124.850 100.980 ;
        RECT 125.040 100.810 125.210 100.980 ;
        RECT 125.400 100.810 125.570 100.980 ;
        RECT 125.760 100.810 125.930 100.980 ;
        RECT 126.120 100.810 126.290 100.980 ;
        RECT 126.480 100.810 126.650 100.980 ;
        RECT 127.085 100.810 127.255 100.980 ;
        RECT 127.445 100.810 127.615 100.980 ;
        RECT 127.805 100.810 127.975 100.980 ;
        RECT 128.165 100.810 128.335 100.980 ;
        RECT 128.525 100.810 128.695 100.980 ;
        RECT 128.885 100.810 129.055 100.980 ;
        RECT 11.120 100.395 11.290 100.565 ;
        RECT 56.250 100.355 56.420 100.525 ;
        RECT 11.120 100.035 11.290 100.205 ;
        RECT 56.935 100.105 57.105 100.275 ;
        RECT 57.295 100.105 57.465 100.275 ;
        RECT 11.120 99.675 11.290 99.845 ;
        RECT 11.120 99.315 11.290 99.485 ;
        RECT 56.935 99.285 86.625 99.815 ;
        RECT 11.725 98.525 41.415 99.055 ;
        RECT 56.330 98.855 56.500 99.025 ;
        RECT 56.330 98.495 56.500 98.665 ;
        RECT 56.330 98.135 56.500 98.305 ;
        RECT 11.685 97.075 51.455 97.965 ;
        RECT 56.330 97.775 56.500 97.945 ;
        RECT 56.330 97.415 56.500 97.585 ;
        RECT 11.120 96.725 11.290 96.895 ;
        RECT 56.935 96.625 86.625 97.155 ;
        RECT 11.120 96.365 11.290 96.535 ;
        RECT 11.120 96.005 11.290 96.175 ;
        RECT 11.120 95.645 11.290 95.815 ;
        RECT 11.120 95.285 11.290 95.455 ;
        RECT 56.895 95.175 96.665 96.065 ;
        RECT 11.120 94.925 11.290 95.095 ;
        RECT 11.120 94.565 11.290 94.735 ;
        RECT 11.120 94.205 11.290 94.375 ;
        RECT 11.120 93.845 11.290 94.015 ;
        RECT 11.120 93.485 11.290 93.655 ;
        RECT 11.120 93.125 11.290 93.295 ;
        RECT 56.330 94.825 56.500 94.995 ;
        RECT 56.330 94.465 56.500 94.635 ;
        RECT 56.330 94.105 56.500 94.275 ;
        RECT 56.330 93.745 56.500 93.915 ;
        RECT 56.330 93.385 56.500 93.555 ;
        RECT 56.330 93.025 56.500 93.195 ;
        RECT 56.330 92.665 56.500 92.835 ;
        RECT 56.330 92.305 56.500 92.475 ;
        RECT 56.330 91.945 56.500 92.115 ;
        RECT 56.330 91.585 56.500 91.755 ;
        RECT 56.330 91.225 56.500 91.395 ;
        RECT 101.515 89.540 101.685 89.710 ;
        RECT 101.875 89.540 102.045 89.710 ;
        RECT 102.235 89.540 102.405 89.710 ;
        RECT 102.595 89.540 102.765 89.710 ;
        RECT 102.955 89.540 103.125 89.710 ;
        RECT 103.315 89.540 103.485 89.710 ;
        RECT 103.675 89.540 103.845 89.710 ;
        RECT 104.035 89.540 104.205 89.710 ;
        RECT 104.395 89.540 104.565 89.710 ;
        RECT 104.755 89.540 104.925 89.710 ;
        RECT 105.115 89.540 105.285 89.710 ;
        RECT 107.705 89.540 107.875 89.710 ;
        RECT 108.065 89.540 108.235 89.710 ;
        RECT 108.425 89.540 108.595 89.710 ;
        RECT 108.785 89.540 108.955 89.710 ;
        RECT 109.145 89.540 109.315 89.710 ;
        RECT 110.645 89.620 110.815 89.790 ;
        RECT 6.190 48.445 6.360 48.615 ;
        RECT 6.190 48.085 6.360 48.255 ;
        RECT 6.650 48.085 7.180 77.775 ;
        RECT 9.310 48.085 9.840 77.775 ;
        RECT 10.400 48.045 11.290 87.815 ;
        RECT 105.465 49.375 106.355 89.145 ;
        RECT 106.915 59.415 107.445 89.105 ;
        RECT 109.575 59.415 110.105 89.105 ;
        RECT 110.395 88.935 110.565 89.105 ;
        RECT 110.395 88.575 110.565 88.745 ;
        RECT 5.940 47.400 6.110 47.570 ;
        RECT 7.440 47.480 7.610 47.650 ;
        RECT 7.800 47.480 7.970 47.650 ;
        RECT 8.160 47.480 8.330 47.650 ;
        RECT 8.520 47.480 8.690 47.650 ;
        RECT 8.880 47.480 9.050 47.650 ;
        RECT 11.470 47.480 11.640 47.650 ;
        RECT 11.830 47.480 12.000 47.650 ;
        RECT 12.190 47.480 12.360 47.650 ;
        RECT 12.550 47.480 12.720 47.650 ;
        RECT 12.910 47.480 13.080 47.650 ;
        RECT 13.270 47.480 13.440 47.650 ;
        RECT 13.630 47.480 13.800 47.650 ;
        RECT 13.990 47.480 14.160 47.650 ;
        RECT 14.350 47.480 14.520 47.650 ;
        RECT 14.710 47.480 14.880 47.650 ;
        RECT 15.070 47.480 15.240 47.650 ;
        RECT 12.240 7.345 12.410 7.515 ;
        RECT 12.240 6.985 12.410 7.155 ;
        RECT 12.700 6.985 13.230 36.675 ;
        RECT 15.360 6.985 15.890 36.675 ;
        RECT 16.450 6.945 17.340 46.715 ;
        RECT 105.465 25.405 105.635 25.575 ;
        RECT 105.465 25.045 105.635 25.215 ;
        RECT 105.465 24.685 105.635 24.855 ;
        RECT 105.465 24.325 105.635 24.495 ;
        RECT 105.465 23.965 105.635 24.135 ;
        RECT 105.465 23.605 105.635 23.775 ;
        RECT 105.465 23.245 105.635 23.415 ;
        RECT 105.465 22.885 105.635 23.055 ;
        RECT 105.465 22.525 105.635 22.695 ;
        RECT 105.465 22.165 105.635 22.335 ;
        RECT 105.465 21.805 105.635 21.975 ;
        RECT 65.300 20.735 105.070 21.625 ;
        RECT 75.340 19.645 105.030 20.175 ;
        RECT 105.465 19.215 105.635 19.385 ;
        RECT 105.465 18.855 105.635 19.025 ;
        RECT 105.465 18.495 105.635 18.665 ;
        RECT 105.465 18.135 105.635 18.305 ;
        RECT 105.465 17.775 105.635 17.945 ;
        RECT 75.340 16.985 105.030 17.515 ;
        RECT 104.500 16.525 104.670 16.695 ;
        RECT 104.860 16.525 105.030 16.695 ;
        RECT 105.545 16.275 105.715 16.445 ;
        RECT 65.270 15.810 65.440 15.980 ;
        RECT 65.270 15.450 65.440 15.620 ;
        RECT 65.270 15.090 65.440 15.260 ;
        RECT 65.270 14.730 65.440 14.900 ;
        RECT 65.270 14.370 65.440 14.540 ;
        RECT 65.270 14.010 65.440 14.180 ;
        RECT 65.270 13.650 65.440 13.820 ;
        RECT 65.270 13.290 65.440 13.460 ;
        RECT 65.270 12.930 65.440 13.100 ;
        RECT 65.270 12.570 65.440 12.740 ;
        RECT 65.270 12.210 65.440 12.380 ;
        RECT 25.105 11.140 64.875 12.030 ;
        RECT 35.145 10.050 64.835 10.580 ;
        RECT 65.270 9.620 65.440 9.790 ;
        RECT 65.270 9.260 65.440 9.430 ;
        RECT 65.270 8.900 65.440 9.070 ;
        RECT 65.270 8.540 65.440 8.710 ;
        RECT 65.270 8.180 65.440 8.350 ;
        RECT 35.145 7.390 64.835 7.920 ;
        RECT 64.305 6.930 64.475 7.100 ;
        RECT 64.665 6.930 64.835 7.100 ;
        RECT 65.350 6.680 65.520 6.850 ;
        RECT 11.990 6.300 12.160 6.470 ;
        RECT 13.490 6.380 13.660 6.550 ;
        RECT 13.850 6.380 14.020 6.550 ;
        RECT 14.210 6.380 14.380 6.550 ;
        RECT 14.570 6.380 14.740 6.550 ;
        RECT 14.930 6.380 15.100 6.550 ;
        RECT 17.520 6.380 17.690 6.550 ;
        RECT 17.880 6.380 18.050 6.550 ;
        RECT 18.240 6.380 18.410 6.550 ;
        RECT 18.600 6.380 18.770 6.550 ;
        RECT 18.960 6.380 19.130 6.550 ;
        RECT 19.320 6.380 19.490 6.550 ;
        RECT 19.680 6.380 19.850 6.550 ;
        RECT 20.040 6.380 20.210 6.550 ;
        RECT 20.400 6.380 20.570 6.550 ;
        RECT 20.760 6.380 20.930 6.550 ;
        RECT 21.120 6.380 21.290 6.550 ;
      LAYER met1 ;
        RECT 9.280 104.185 56.675 106.365 ;
        RECT 102.030 105.085 103.225 105.455 ;
        RECT 2.000 102.000 11.465 104.185 ;
        RECT 2.000 47.825 4.180 102.000 ;
        RECT 11.645 101.745 12.335 102.205 ;
        RECT 11.645 101.155 41.475 101.745 ;
        RECT 6.620 48.695 7.210 77.835 ;
        RECT 6.160 48.005 7.210 48.695 ;
        RECT 9.280 47.985 11.320 100.985 ;
        RECT 54.490 100.100 56.675 104.185 ;
        RECT 56.855 99.845 57.545 100.305 ;
        RECT 56.855 99.255 86.685 99.845 ;
        RECT 11.625 97.045 56.530 99.085 ;
        RECT 102.855 97.185 103.225 105.085 ;
        RECT 55.955 91.165 56.530 97.045 ;
        RECT 56.835 95.145 103.225 97.185 ;
        RECT 101.455 90.085 102.855 95.145 ;
        RECT 109.625 91.550 111.810 103.560 ;
        RECT 112.110 100.770 114.295 104.830 ;
        RECT 114.595 100.770 116.780 106.100 ;
        RECT 117.080 100.770 119.265 107.370 ;
        RECT 119.565 100.770 121.750 107.370 ;
        RECT 122.050 100.770 124.235 106.100 ;
        RECT 124.535 100.770 126.720 104.830 ;
        RECT 127.020 100.770 129.205 103.560 ;
        RECT 101.455 89.510 109.375 90.085 ;
        RECT 109.625 89.365 114.820 91.550 ;
        RECT 2.000 45.640 6.365 47.825 ;
        RECT 7.380 45.640 17.370 47.680 ;
        RECT 4.180 6.725 6.365 45.640 ;
        RECT 12.670 7.595 13.260 36.735 ;
        RECT 12.210 6.905 13.260 7.595 ;
        RECT 15.330 6.885 17.370 45.640 ;
        RECT 65.240 19.615 105.130 21.655 ;
        RECT 25.045 10.020 64.935 12.060 ;
        RECT 4.180 4.540 12.415 6.725 ;
        RECT 25.045 6.580 27.085 10.020 ;
        RECT 65.240 8.120 67.280 19.615 ;
        RECT 105.435 17.715 107.475 89.205 ;
        RECT 109.545 88.495 110.595 89.185 ;
        RECT 109.545 59.355 110.135 88.495 ;
        RECT 75.280 16.955 105.110 17.545 ;
        RECT 104.420 16.495 105.110 16.955 ;
        RECT 105.290 16.695 105.970 16.700 ;
        RECT 112.635 16.695 114.820 89.365 ;
        RECT 105.290 14.515 114.820 16.695 ;
        RECT 35.085 7.360 64.915 7.950 ;
        RECT 64.225 6.900 64.915 7.360 ;
        RECT 105.290 7.105 107.475 14.515 ;
        RECT 13.430 5.080 27.085 6.580 ;
        RECT 65.095 4.920 107.475 7.105 ;
        RECT 65.095 4.540 67.280 4.920 ;
        RECT 10.230 2.360 67.280 4.540 ;
  END
END tt_um_wulf_8bit_vco
END LIBRARY

