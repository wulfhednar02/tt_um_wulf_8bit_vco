VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO (UNNAMED)
  CLASS BLOCK ;
  FOREIGN (UNNAMED) ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.005 BY 0.005 ;
END (UNNAMED)
END LIBRARY

